--
--Written by GowinSynthesis
--Product Version "V1.9.8.11 Education"
--Wed Jul 26 12:23:12 2023

--Source file index table:
--file0 "\C:/Gowin/Gowin_V1.9.8.11_Education/IDE/ipcore/DVI_TX/data/dvi_tx_top.v"
--file1 "\C:/Gowin/Gowin_V1.9.8.11_Education/IDE/ipcore/DVI_TX/data/rgb2dvi.vp"
`protect begin_protected
`protect version="2.2"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.2"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2022-10",key_method="rsa"
`protect key_block
TCCHqPJOsRhi9Y28WJTbQjMKVAota+A0AlmpZEyGKv2zZke15ulZ1gj+0iiUIpu/oR3BTGsb5xqh
0aElaePZMEBTWcoz6qEE1ryc0Y27zpUaMVmcsUT4exqSdYf2soS5rFFqFiQk8MZdBV4jyfKkhzda
UL6Twq9o+w44Bi+8pwmbXEyuG5etlnLBocLawC9V2W2uhYFhG/Oeq0LIWqUyu4vJynO603yLtGHW
NhCx6+/HyfYHjc2zjdNGG3u2+Pm226UtUO3/vm0DYaGEpIiQ++HuNuXVZ4AMrYFQ77TFxVVc3O9T
mejDwB2J+3Uglpuca0UOsTSu4GG5FCcuruLMFA==

`protect encoding=(enctype="base64", line_length=76, bytes=67248)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cbc"
`protect data_block
49458GRtkhai5dpzK6i4o51ub3JNQV8Y0e32O4i2jiw2/a/znbKtH3fV4IbwBqVuRo0KkrI06HC+
kL7kS5prbIIp7GwOtePr/oJskglJUVohI1R4+wjO+EoxTg1akul+E3LnfpUMloXL+nmDL61yRzp/
S2QWCg+1xpsRgaLi9ICHSVPoEQ91Y7O54yjHTFNLmmdfOlZT4b6udXbPanevOCvHXP1FFlt11ZKx
AOnK2dnt7V6ECnI0w+XeyJMup1QNJhbY+h+vJb2++UpVczbykBsR9nZCHeuN/NBVT78WWxo1/VoL
JgcX0IzwNmbN545jKB7/KE50e5CKEecyKh5CQhsVdZOFKd4aWSTuNJa8SrLGDumeE0ZQlMOPZZCZ
yxzNOQyKkAxZLwTrloN08F7UkSae7/oO8p40xWe6UKlvwcTOG3hbm6GJN9RGD8i1aJG27oYs+Ndq
/KP5d28+kfQKbkRMlZsXw5mia36w02Ymli7fsk2PYRaGNO4ACMIVJWn6tcuFEhXQ0YIF82ErZMHV
dkClpnmkfLbYpz2AxATd/hWGB7hchjEp/v/zV1/kjXriPU9ac1MTEDfZ/QZl4wO9wnXqneqohCUv
zE/eLE7XDcthS8ONr20+UXsGYa5/hMXRm091M+5WOQE72GWXu4KtNs28mvwo3knnwRIUUrrvaZJQ
oVe4Ra99P+gs3yPuTNEhs9iTnvN5BuCv3eXQ1tuzRwB6KbYLnUb2tXoJMW3R1gPt4MSsrQ+/lxG+
yBAi5i7UWqId1Pp+Wao0qivDfeCxN1roz8X53g/i8AXvuVBqTftdmuPSKylhNiSWVQhlSKCpyNPy
FxOzh7e4HXrUpc8w5ILfAjv2lJ8irhn8FfoUJkHcLOSBV8ynpM2QR22gT4Ia97BecXwWSTZ01VC5
nYB1WZvogCu1vgubAJ1lWVXzpQtoOlo106G9/B4QdgTuPiP5Dlgn+8Gde1/yTvuFYH7ROmHgR6QW
ndnfwm6dfKOU3qC7D/nkjbmpHWKvfZhTnrGLdChShKR3GpyEnCZ0RxXRoxDJ1ahRkJzbu7dFzJB0
2kMOKVPPiuhCfD1qibelxwUPgm7VVWjG7RI6dIsLjZ82EZjoo/B4y+ab8p9wYrnE9QUGKXdOxH/B
fJ1liuq8J/nV/8zuFVtdMniC62zRj5RtnEcho9H8xRmHLBEvoFErLVbXji9wcKeva2Gz43s8W2Lt
UPmT4cMyt24DYu/aBFw7HiWBtNjDqI4rE7QS5yj5Xw5TBBm0ba9Tvt9utG6P7cG42eYcJFFuDlZN
JQ1At8YHhu+d8jTw6vJltDDShrGANlJASGHlkAPuVkdw3Km7FFEX4oVDTwmWYc/XSzbJ6D7c5ANb
MUScQUGRg8Z3UNENsjf2wN6qZHkjiSgpcHY021I+/zgHHA52BmflKxJXyPYTOnfgslTRraMYb3z1
A+6tCHoHTyDEnXzJQKXaU8lhs4vNoE442S3CJs6TqyAGMOOdQgRry1XEEcFxKCbavu4fVmnWres2
a3nIzrCF33BFcK+n9jY70mgKb0EuEL+TXMD75LqgHAmB4+xEzvujA/1TnxuV67jmnQbfMoI0kYU1
C3ouwUI80o4tjyS1qAEyPX80e6oiO/HKDsBaBF/nhCAaNin+gvZum437eTejYIhG+yByC5Natfcu
Sc84ygcOKRhzxDU1SfpzjdSf7BB8PxcQJEwbdF3k5oUST4gMizo+RjDLUTsPTqzEs+jQJctOW9Xn
5+ggPjK2ZMnTWlZPtm+6lgoOjPM7VM2ol16NvUHewXqYPyV3XKR99b44HtrzJ0jCUtCT6aVYf9jz
GHGU2xwcEJlA3h1wTASPHDJTMjNU4zd5jFZqLHN1NdHd+nO+O0TjWW6hSb1Fv151PbG7qimXvSf9
4oWQtUWePkuXvRbA7v//uke+2F4sbOzLKP7Y6TrGLdW82ppd6vsy6Hx20WRaOLqVK886w+QgNPmr
iLSbux7TAsFz98Zvn2TcL0GOfa/hlCP3Mc1BDDVc0EzrmlbQnJqUrBXL5Mf5mFOhmQDcGzOspaNk
zc3kJTYaRLwPEnAd/VTr2yzXQoQ+i5/HTqIBftfi0J0/SxEmjeHZefzeVwHOTzDrCQiMOmxaqNBa
zNZ968Dg8Ol4U+DmFG7Hgaxi6nhNIu8kYkrs5KF5kK4WxcgqsxFMf369VviNPafOK6PZi2BxDwy2
wMlwwhN73GEzLtWXjAO8rQXiiqd5j43IXe3SwvT4HdMDWvkuA84N6PiX+tiI3g2ikCidcYAHV2sd
As6sDeGBU0WclXlXuj2GTzYXW0aml4eQ6T8AmaPScsdAiFAn69chaqxdaKCfVrtyQSPfc2VFfN0y
kKpcK5dQOEBYTeNAVgmnp5qi0F+6zESBBAmhCSdYsxq6uXhxduZCTQQXwES079Gu71qikwLd5g/C
osc7LpbYcUdMgO/psID6vDJ+RwlRsSBI5onqPqL4+4MWMVIgkGDPPurO1CKdfhRkN2mnODbR/QMD
UJ++m1B/3Bj67EvoVVtkhBZ6kmuvo2Rj8sASGH68tLK2TzVQXhPHLBKS9U77sFhzTQyguMlLRBA9
yLwBs1ij7KrM78mgk/6VUbyYmsxJnyOoRAYwj5b2QnoTuCrINU6lE4jcchesB7NrDXjLyxWc3YiB
iV1E380CceRQR0hhdF7O34aDf4vIEgSlt6chnbDlMrn+ByLK8MugVM4rRJtQkNJtJ/ECE3y2Ib32
4NHXoqIhbwAl3PkI2nz7tNv+LNtIIApe4mr7XPbGVPOTGPMy8hxNpieZG662bayhu5+sP+SDa5EY
W9B2nRgflfuhxFdgO3Ij4M2k/BTasgVT5p2exEtm8lQwBiSBNnfSMZiGW9rplMdKxLW7lylmPxJA
OJgwJnf9jEheXfdiI0ceXX8iOgrOmCL2w2ZO1ea7FeRe1X9A7J2yrtAvHMHkctO+L9NG+Q/HuBDc
egNxxeBspj4yThRqO1QjKhAnjb8rHlu0l0d6TuUnVK/qvWAItE3ao+uWl+ENOqRyS+QbSdcQouT1
YCAML95/2kt1VuwVIayqkHw2rHmCgAW+Cs2E0ZiLmlNc6b9IHFulsW2IrSexk0mh1Z04VGXenIkJ
Jz9Y2tgCaaxU35drctz5Hqk3TR0+MDz13ZDiAUgd6LQjINKQGzVwj8S/u6fbc2npIfCsNLHKpiOt
vOufievFhJo86S3CUYdXprGPXio0RkdW4jF4NYfuGn985IoIbQ+nm4cW0NbQYSmNQQSHx8jsGbpV
z1HODuy+2ETqH9m/SrRUzE/4e0/uXTPKByfvXTMmtz2RKbyzWkxOyn/KPA4uULnuWDO3Iyt5ga5+
L6AOHcxLJ1pwVvXQ9MbTzmW5NX3fn21RB5l1zh4AQ7NOiISpt1sxNU5MFxkfNfOxETHoF3zsngUT
Rov+vuqKp42G/caV8MBkBuyM5bRfARKGxitU4YJJz+ZGyDI7v4ECydjP8WWXpb+mV7HgCjHsRQ8h
nlbmjkWTqRRpUAcI9LYIF7j9w/UM2dKzWdxKLyThSE1HbsjuMfwrGJc8f7itcFmcVSYQR2NGPxuw
bv6wgpvNl8avkrHxkyZo9j9B7b2VqEZnmjY1dIPZBUWNjjZExLsgN5oxR/dkDP5Ixl7bc9wtmT5D
wOOwt5nnGkM/SMfURkSmTWd37ZttUKR0p5D4JF3UDx15v4a+5rivwdvET1M0+Lb7BD+V9tbKdFsp
FAMR1VrvLsphO3uAyvtJsrSYeB/kvVQSqxdPttLsKzVDycDMyrrEX5CPrV+sYA7MFpOkl2nkrkTS
V7hzCqELQv+GB/tHZcP2J5w9MNtKryxRhv54qgTX4/LSiClvnRj6Gt/pcyjmbA+D0G+nx21OAWr0
yFR0LoI6Ux5xdEdusE9o4nfeh4aOTFTnoIf1xVMKzBQLrZZvO6UZ53S+2BHEnWd7ofGKXJCcsQOj
uwTHala1ewHHolSC9zKkHlHAV8BpPjKo2vMWkkeToy1/6MT+2EUUeVQq0TDtSAWgdGcmulY0hXWj
Zry1r4mPOjQ6VVEknZ1KGS/O1sT1LKq3r2lWHRHp8dZGbqjdOJx/aqn5S8Xq+Uf7ODtML2ftJGZ2
kZ4DbnvLnypGazMRKIeR37sJ8UbiztHTTsotz7vw3uv2n7PNxPX2rsi1XukQE1B2d+p8hDoQmZPZ
rsio0BYKea66GbeYsGJ/HdvIocVHWqEIULEShdRnbcAJOJomxkrq13XqVieybZiZ7nDE5DHyBYYs
szcq4cKEmwnwFTIdc79qXLVbveZDw5wPLjdCZUcEvU+DevfPsSYLOL1h0A0ELI5CYtzccTarxMiB
nbLixZ6QwC0z2HTiXqcOrE2dV8MycH7TwAlTQI3SKtXXcafwiekVWszx1i+ZJ6GPjwQgO8nVnuGL
R/kl2ZceIWlYmdlAWYFgfyuBwHPXC9bftH1Xs3XiRKcQ3BHN3csKu2t5rPGlUggJ+laTuZzbu+LG
oGPo6dfvYuC3NlHug8ALAuW4B1A7yX8bgR4XrgOH4fqYmpu1FELJkrGbNJr5XDEx+jCJ13PFgeYm
pb9pamRx5vys3wZ2S8a7Gcw5sAlBHrjKhaLNSX/vZu8GYJbyiJRJy6SFO71rQrOS8zhCdrB0FxkV
7d7yyH8wUA/eeotqrM/N+tWY0Bisoja6cjpHN9PtFjUQKRF3NXVK8jdO5hKOb0kWSUZ5NDWteqme
kB3U/7oN9FTLbbtTBlL0GRyiR4wlxyhtknpvjHTz1uqo6/GjvLG7rtOU1FQMu5rWvVjVQN416VFR
5UtlyazMNGwzJ4q/0abaZXUtV8MgmF7vNaOFprKoPDngTMZv5g5k5ofPQtp1KmIq7L3V2P64yF8D
66MnyjglOM0W0kj9OzEaQ0JVMLcoGOE4EUN5zozo0mKysM3vbxUbIoDKU5G+8skYZam25A0lSo2y
MQJvL0JxdKACSpGP7cHS0pu0nStU3M0uwrfV+dLAyyRRn/EmuGcyWLTVY00rqun8MW113BocpGK4
wmXsMtW98gNxY+vz0HuuXaCGzMH394M1FmB4SOI2PxKTpyTpCSAMaWgoVt4cDWyP7cmF9dReDLEt
9XJOTmBMw7cQ86qfBB7bngQHHlDgoZIrq9RVR76hh1LccbOaLTIF072rTIsMabk9PL86LLF+Tk2i
HXSNT0Ymd53llbAENmvdSJvthLDql7HZZgVDPnJkUtFDkZkFoQsVrJr2kSk73/B0rhpCvvlBQSsW
T3GJ+ZK/eFbRDufvCPHV+O//fPMTPl/XDjkiQJrjZvdeFQCMgOie/ol3dDwXntNMJxCChcHoRSii
I0V07yCQVznnPFIKRnGn5nkegZbtEqNne4sALtex6HiSCDNObupC9+mLxL0jEOKf2GBRQ/dJBh9d
BfysSRgExunJodtRJkWYnyo/mJHAXtV4fw48FD0uVG2Pe+gHuvCfeIoYMqOW8b2hNA+fUYaLycos
irDkamMiFeIw9cznNzHxvFOTH+deb+tOsczec26y0olNv5BiOQedst1iBy4wIN0x4UwgU8UPnCCI
RT3iJqehQ4avNCBagK1bG7OBY/T0ypG+KHTG8Hm6V9E8JSvAfxmjEO4tQCgiJOEUx5Y6mjNQpPtr
68Fe8AAr3fK1VCRVLcFHq+crMz1YfFHEc/rD41fUY7aEj5FnswETAY14W2eMbQ2K9eZhswYSZdQl
TUpBxXjcl5oxtqaHs7xUn4xdZ5+tYEHBQm1/MJHQUcFuHvV3XAPVgZM4WhULEK5vRWNfsMq8tuXB
t6kXMUjLQdiFYtwlgpa7Q9/M3PXMwDTwYX1sCrI1hUgfSjPZTboOvoUv1UGjnXJtTtkZic12zMBp
TJNT6pATbxCUVBfN9IKqb6kvZ4U8C2aw2yf+chNWa94OuRMfftulgal2iI75GgX0hVJ1SR3f8rOo
F51DN0HW640lw3BpdXltDilGbV9jUf7eADWujrcX7TdYxUvLZ7yipW2YoU+htcS0S9B32Yl8a44C
QYKnesjmbcW7ogSeVrjiNoOfVG1mK48LwfQcAGG8Lg41UTFCvIwqPTDaEoUo2PpeBk+YMKHay8Nv
d/k2RGulj5lAViTzyW2b668re4Zz2jb5M8AbpFfVopnr2ueaAgivpUO4kSQl1LthHC4D6f7UmUyl
sxSRnyBcBOI7+IeGxgjUpX0PphzBIDnhdBOWXpgBj9TAKUsdemEkMf17F+fHNOIdd2CWAm4TZR/M
TnbQkgkZ6ZOxneMDx4khGOqc0lKysxSNLnek6H7mvcTgc3yRjz42BuELMgncUUKIxIqf0xeh2vS/
Zvo1TblW8LSDouUnGh1aT4Cm3OdU5NFKaxfCDDdxkPoD5mJfo6j24nQTwqckKeVlTaLCvcAsb8E7
ILkd3hjkcUPqkvm5viSjOnB1MdVs8ibI/3hLS25+NHlbvFV8kUDLMVJH1tL9WPrNBMxUBoK2tdEb
WjthpXDFNa4ldjvOuSNPl3d3Ax7cHS7AUyuf7fExMuluCprR8yCLR0+4O6kPx4M3uKgrS/VsQwNQ
VKb1R6x4NOWgWb7q3hMYZUgU+yTCmQ8Hw53aWoKeOp3aEU0gY8webZy62RVQn8/3t50aT7/X1Ur+
OkobpmuSoG96yZHPavXJXrGw8nwUzQ2Hvt+OUYbCQaEiI0oONoJD1uFt0tIwN1KK0kQrm+Bmu1uB
s9cuzsMiogmdgH7rNhMj+NAAs1RaM7Pooc3nthrfBcQC5bc0FkMh0B+quMlGbSbA942Hm6uVBtr2
BRq7YjqgqX6K1dEHsKUVhLgo2pl7+428xeXzdx6AJMtzALGcmNIQ9ijyP1qQwamOgqg4shNdo0Do
5/CNN9w6gJtoSuYyAiha4m4gUL7A9VwSrjde38q5rO7oQAUNKifKBGy7/LUJ/ur5PwLeiJ2Zvlge
xYhSpaDKS7IqTDdR8io+K5M/zrBslgPJMOfE9UyzF3mVEaBcbMXkw3vHPV9Zrb7oTC8ALRB/0bmd
UW8qcFVgtBWsf9GIRTN7xgj8Yr8kYROUYTvmC5Xgpg/oEW8Plk/lszY2oWFom0Ukr8YFrjJLJpEj
kQkU3hu1Zi+TcRLeLF+Ckn3OgKBzM+vN5m4X/R5TyRtrZlfMleQ0kuhJSqBHXWhg/0bt72fBaE9L
ddj1Cxb1/bjovnEQc6ycQ8e6XUZujH7diYEhy7kl1yC9D+AkiCySnP/qzJtAWPU6PV6Vw21vnRxh
ZE9CC5ls13hz5G6jp+UVQwZ8XYmH8BXxXIwbNTwiKu1DvRlnhIGfKDHf0co0DVrDYWQ0DMoa5Iva
bCuNNGxhQ4wEyTNcg9ul9mk8z31vG95y0szchbVpa8mgrcr4ivQAkU5Rx4yFTTg0UB6iPcm5JcDF
yFotZtGpnUWyTe+59N3KbzN0aH5DKDadMtH7v7B/FrzB95tnj5dYncQkZvDuydEPi0kz+lSgTeg4
KrQzG8d0mpCYwGfzNWhz2RGcDPBQ2o869Co2Gvqzk93og7cw7f1LZ9e9prjK4ibtQIkWGkhG3or6
IpJEdjZBjGE7JGplvmPMvLfyVCJZjU9tM/qGlTcwZJpBXei/gp3yIpLc/VCvVJMEQhhVUZagJfGu
GH6uqhoh0CWRBlyR9ydRVdWKiyJsMVXReX69s+o1IJDQO+waA8vSAHFEGh36CtY9jPPrmUbeIfYA
9PD2OW4CvLV5xI+0OiYqTVBISDnDZYcNa7K5kmcSsWPSzw8B4YgtY7epHfrE6zaq5nYAqFRJq4Aa
RHFp1cpqFXCjaId8xTdJfxmcAUm/0tMFokwOVbcf27RhN0pS28LpaW/qvnhR0FY+QCFCOZy9Pinf
ohadvgOytG/tESObVCGSAWyPMbNVHj9E+zsxWOMYepC84XK1Iv9rx6AKeX6k199d7NYxPlzsYXUA
xCrywPKpo/7/NNlaBPC8BG5HffVTk+UjP0gq3jAa+aaR2XTAUEKdZbcKH97eNzFiG1NmrcM4I+vf
jJbYAzjHidQYq/G6h1YdjJCd75XnUxVZZI3zAKKMrSW0+Tc+eaGQzgJ5LI2lcZFhgjEl7xcelpCR
xkh80LWvkJTUmkd1rQgDivwDBTnbsabdFgx5keJeFXijSUPU74rixfrURimAxQnK/PimTU4Q0e7z
K+XGKlmgyrPpVE9tCZbjkp4telEQbtJI/xVJ3UiBBHZrK4tfBMqhnmmn03XllJherzKRF6bTXJfj
tBW6kXGdpFEp+25+vHMnSOd/ynocvYgv5spv/RjDivGWDGMWLhDf4hWeZyiGvMeg+YUllcCbtLT+
LJ09k6OKtoircb0GkngFA0uqcVOB0uzxJKVwPg7gSgR8A3TErCzK1ekjQ5WXP4TS55/naVrW00d1
I6V3dbkcLFOw8Hq8cCSKyPi6c94jmDRmTzlOX5tsSdP93aHE60Uae/gD3E/gN+JsVntIl0qyOxpJ
4Z6UrTP80CBc9g7+EZPBPCnpfS+rP3UFKUk8CuQyt8lpwW1Z6CkFhkYncG+JcCSvLIX0M19hezTs
mar2PzyFR3VL86P6IaDPne6Gwww625ygTj9iNPbaCSM1ZCE1qatdtNHhnmn52cv0BUkiaQ9FKZXV
pfdJiLtBNrqkmCEqy9rlMhkdTwAVtfevQ9RkpkUco+fwS2n8zJ7NgK5EdxEpTyTXIYvR5fMUgjHd
PU7V0npAHD9if7twUPNOLmG5Zo95eQ+MORw8Y6mD3FeLWdITQXGJ1pxVp1UZbPn5p7e00VgzeIbB
ThcoXFwwFSJbolucxphfUsZ1P4mU6mhaYncRJrwxQSAqBQnSKZ5qjy3G385J4RTe+AKtldUgv8ej
tarVoQ2dlSU1cce78J8nb5BqjwqbnahzM8cdiUFe9bq3mJHX5KQw/cg/04esmsB63325mAOM+ISq
IXrusHSq82KHk/2c7jCvGR459ksfrL3uo077emKYAiIeTRBxe8h5fZJJfSj1m/7FOl06oegqPevQ
j0lw4Tk59T4p26OgDYCxV/NR9L9IrDSLgR5cUCuZinFpNTpgx7QVWU84vpZHdNn4lI0g5x5K5yEA
z+b5MSDcKrEk9zRxUD+pN6pNmA2xgYecrZt3j6PNj414pL6s/q8XQVE7pEl9afuUMDtyLBrlMFFO
0xS8XB0Jrb5zoWz3EE6GpYEkKgoChzeH6mt9MREj+A5KhWQhQBEIjJNghWhT52voBrtHoNWBRwFG
2sR88CoggEaHHnb5HkcEE+nSdNGba3b+Q8/R+Jur0yYYLzRQW64Hf6QSn75UW7prx4YrsPi2RSHB
pfK5LCK2i7WR7iBKdMQGF7dKhCAvP/mKHOPUGmJZ1GxZmHgCIG9gXzpVnB/jMbevyagNijGRcq+P
Kh+F1lI4Wu5CwGBRIlDf+Pebmg+HsqrmNuiBjwcDv29y5fBfWX/SylCzMERRxnXVloBUQe1D3aXF
02qT2Z3bLEtukUF8Aglp1M7gvvNocjii8ZnW0Ri+lRJIGw35x3i3wsIDSiDlTGs5ofKnhd0/iyI+
HJp0IzGFBhSXUT8XHdipKGFwwZyNECFPRO9Ac9P+Xv2kjn29NJZ8WjeAi48gw1141UrI5KkcYYyL
E8fMzQrW8f3VWaYHFLnaS99l2G2e4m4ldj5zTYv7+ecXWBDXbgxJFI84Ic1ltlHaqhEbudZWAH0T
cP18cPZILiLSgsMygTcS55fGmawk5VEzUayZYx0g511mwl89ysNbyYjspZF4oW9tMQ22JYTUUUvs
5fHise3uvtOOmpi564YPV/BqMVDovh8TIGaXPhYiGnf2qT7YFMchSsuptoCf4ra9N8nTUX8Dt+kH
K8Sg0XRFyqOzOBWYhh6Hs4fSA/pJj2kbK1110uApoWvVKH+h7myWS+BS+K2do8dPKIGLNTYqn7F7
Vv40/J2K8uncsSxeDbuIiV0D6m4AJo6dG6uogYGXBmSdun3aP15V7vQYrzmc8QukIDcgxcHiKYPg
tzAc6P2xstQ+o1On9obV1QFpdfKNpU6QAE78QI4LXqZ8cYTzy2DYyPdxq+Ti0IH/ndkgpJOVvHkU
zHElyDA4+tyhM1PsTYSYaEjb3racNdyDmoQcsIPjr3Zn0q8qv9P3RWJ51aKGZAmKvNhfuIfZEno6
a05DHgKk+j6K0gZ69X9duxkHN0GDe55JzL8ChV4551s3JcF0jA2BEuZW2ZWNEQ9DoHPHgStY+XHD
dGBGgjdjVWhZeRkvBfRpEVl16nvVuYcnm7pHyy31vsEoy84uJRUeTL/2QwAsrai/4b+v23BDWaPR
VWDP8at3JT/Dzhp/kWFFggkGhavpngHqbADg1AHSnrFqgGuj7VSYWE+nkaUF+0QpOgcLA1tLjpz6
1c6PH5B5I6ejADxTs9qXjRw5AXrAlLivVhsP6xuoDUVqD65EF3auXi0/eYU3LV4ZoRF3KMWe59bz
g2PE5WKr7tIZDEPpTonvsVpRgwt7Twmjb6spcI6YBFML25sz41nG3uGDZO26lhszvp6ya3gV/Osz
is3Gx3ORLV/jKVksWu9ZNB1b760hX8KFjKZ7PQbPyYm/SVznSDFF3zNXWSgfKq24fCNRmLbMCerm
nT9WrfbjK2Vk2pi4yidjDYv6Mdds29bf+GGXMB6J3LHtXglxR9bg82ExCfJbwMKldwE2mgX36NgY
x0inT1/pQ36lwGEis1b5cEZlFAAp7JPHROvED8EUZIi6Q0D0Fq2bo3gTD9/63bbdVASBCjPIKHdd
pKgxBG3hg3c/i0tYJ8nqrxPSUndBcjL5i0f9VPfKcMtW3SPV3lC8dWktRnHY4MbB/x2EHkgzECxU
CfK9zATl6W9tH4KFMX9iUqnWIXOXJfJnAY9uRcRgZjbSVs8cjD2s/6pI8K+1Yz5nagZlSQJZI6Fk
B+8t5eRduPIJ0aRLnxBlPvJ9ZMgKZLo7qXU/0wTmkmazzju6FJqALTsBl8D+HH1vH75+lYY+8f8n
325vi3O0v6Cqyt0HrgNhDqQj6eKhM/gBX5/lcIv1Vc+4EFHqzGK+geew4EvNKHxcvMSFUJHQcQ8/
dCCrTazpCXBPk70PA1HFKC4H0cvYh1aJ+KB7b09ZBzvjnkqSa7rzGhd21ZQ2npBo8fY7o6amYpZk
EpEUZRrK6VKuInluwERKK8ZgqmEmJtPuwY2xZLxmaaoFYiA4ev93G5V+YLtP4YRHrYM0/Xg4okkE
bhN465IOqLqxGP9ZnVYFSK/MdIn/8Jm/bwUCR996cz5E/j/n1aFjNQJ0/3cWv7QtX/lHtSu51mhP
WSIiW6PsPWRoWxyVpQHcvgb+Riav02OjRL7W3ZzvrAN3MPfyaNh2ejdx5NzEVCmJYHtV78t/T+n1
0SQ4PjeFWN1r06TxuD3dZ4P7JQIndq34w+L1JqzXQEs7ld71+q//ZyBNj8bRqUq0bQFuhDBiFBTV
HcqaGZZeymKipT//Mi0Cihq5WwM/pdTewD5uXQc9RkZTZiGNJcclPtorcbgCnkAQ6DyS1y27FFcF
PdUsK7e0rZdEaA9nI81d/iPaWx5CHsaDIY2wfyTOJMYkIYN8sAhyT3hptytD0DCQdgje+WkN5tgp
fCctIgnbK/mXOTXoEor3yI48hHRzJE2zdc0LByDDG19aOynVA4jTXjrEQxwlPiL1R8KBCYxSERPG
y8ja9P9x4ifaHYX05T4GcDjXcW66ltRWkyZ0vAEP8RJmSMYBgGXTWcOd153PtYtCKAfEngq6nFFF
a5qmFElq4BiBcwLnqg4pITNlXekXpZcpD24Qg11QS9T/MD8YMNT0PDzn0ad5MsrxfkiPIrXbKLLm
/QwoXENwovwOezJ540cXgOlRKyQdf7ZG9deZ5Dl0s0Le/4sVLNw9y533GWuY5UGGrFDKp8EMws38
RgdRfa1j3AeEGPOOTSPL+85CvFwaxpTyvSQmegblBGCgIjyrRSm87ByiWZYuWfM+TFA/OZVd7HCe
oVgeqnQgZatfwga+i0GXZJcphHGQC8FcXAlT+5uaToEBTD2pmLGOfBm3YkQY0q4U5oCoRCG4ixDB
eVmf2bV9TNm/UTWUADgJYEdq2akKh7fXzZhU+3bZsiaS01pWNkSkMt7iFcHRzITgoP/jzCmUIYYy
vXxFodSlc87ualBNbKLYHkWMTQCsv2lr3SLDtcVjfzmm7Qp+7QAHGeR8lAiSk9WOGLMp/n+puVuu
OWFT828qluthun7PDWfNs1PzgslTnf8X0hvJwuln2HaH7sAtHSmPp6ir8BXfIHaRVbrjUCRoFxO1
V9tUAsuw8HENDVCe7emfHDONpjaCvnoWBLPB4Z2VaF7ta1XQhtmiaPByeCIIBacsova0kGw9uUY1
OX8BCOaQvQz4FlkCJQycNjlyl4NjclROsR9UR2drFhGhhv5edj+ovnYdSojnw0ScwKLjm8xsumhu
Re0bw1rF+CabeLdwgIEtqLbowGDqLUeLBb5z0DBoGmHFoHRln68eLWuExsp86pA3oWCYgz06FBnl
KGTsHyYLvTPxKKhjIuQbaCQEya98rLk6DdGQqAKiMZEQAA88KFX547NhgXvxXufOyD1KNrPg9J0I
MMvYoeA2Q40kN4meHB4F8NsWjfRz+HU1dVpvbq6PpwE9guoBes5S2VHDeTdjgOHQaDorUojfKhP+
DGB9bZSEUrjhdZ75363B4CADXU90nWGiS0BxVpr59lnZca+YnyG31vMgnVwF1hLjsuYT1IicI3+v
pJzE4ncejNozqa1i4ulBHUb1eHCQDWHGakuFX8ZhZ1QfG5dTKimIunYZ9JLBHUCBlCvL8Qq9ZSpu
wHs2Tt4hvUxJJxz8HavL+qwaok+IM0Yg0cK6Lrx9hhP22QK46eg7hhNDH1Vgf+w3FB8XGcD+MlrF
ORmubGDDYEizqsTmTtJBt+e0JLzExBSmj9nG/tZzGVIEU+pFf4p2ijO2Q7zNp1cFfTs0AAAp4YuA
/hYYFkzUFJPJ2xCNUw2Cr8PuH8ElqdOaHzeehhwt9sWUKR4IGtvAsf2Y0X0rbjTNwJD3BbmTq9SU
dCo+pDiXFkjEy52KBPIKa2lU6RFVUHcVAbs6VmIY8llNdV96X+3DdC5hZjYUJPcSFZxJB1TA5wG5
bmI6kRyhf8KXV/ssVY5anL5Ehtd9PeU/veebDtnhFtfYyZS0I2P2g1MRyh5h8pjXdQ5YZ+SXi5YV
7VnsMChhz2M9kt5VjurJBWBM3NSD88qU4PXwJPCeJ14nhMDZ308m9waHPR0kUrjg5O4z/WlugHkq
fNcU+aXwWwHeO8S7HlVD64MrOtBWMyJF7QqbfAHn3M0kqdyBhp28qsEBhKS6sddKp5ETcFVttgQj
uya+ud7VS7aLWzZUTFfWStKhRO8Av0DrhrhlOD1gMYcXWEyACjPvUV14QhoNe+dqX7k2EvFPEa+9
pW5Ycoq+35kIFIxGIZof+wF0HkhJ89zGJ9Xo2R92g4i+Cquo1hqsf3eBNqdAIdqgxtbyuVCd02jP
qtKbOKD0x8BVfFmR5B5dKOzqiOEaitJ5yoE/G9bbCbQzMte+dmI6nNOtx+DOYKJaNNYwqaWifrsO
wnukqMPVUwVePBlKdW4vE04L8H88kAheMbYFRvIAiaNfbVd4SfI+v7MJP0wC+W9tNgTsE/VTdo1J
1+/pQv8FUP2uJtP23qu+11VGQIgCssHvnnlz1dSclw7tfrWocmHLUPey5FMHgIV2yo6mx++/qyav
cOjiagfWILJQOPIltolxJjPXYIfduCQyAcfEJxRn09HxsOHQQ1QTCRXutEjN8gg5yqfcwL+cdc2o
BZMCda6xYBGdjMv28Z9IdfPgNjiphY8HhDvELpIu18387o5HZbFXgbnZYwe09ssmkI6dzC3G/Yg5
MVLKgCr3jPBsh9aTY67cgvOLrMslK0+M121PQ4FUGq0d8fsXrPP4UQ4ApIORoRBMmWVZx4QRgCc5
lZaHvQ0iS03yEgfOTgBEM0+xb3Zdn1aLkIhbOCWk83AqAbUHWH/0d3V2PSJ7U/FpnWsXIaQlCBuX
gxTMXWMBD4boRHPUJqGThj9iqYDC/8mpKaRrekhtBni5KSGTxAqTajm2f5a3Ze7W5g0K1wlx14VP
WncpJv+p7Suad2OsuBhoAISyzk/i/saCDvpwlhLmC8Yo+uS1mXQyksndfezeN7hDbnlJHvh58gvh
pu6PJhQRuiL5QJqqeVpkGc78ADTjOrbGTWeoSBRVWAduoa0LT2r3b+un5GDUjEqY4USU4UfIqZDw
zBp7AKNKH6sFhHlt9zocDm7nPLjWNAIORqJ0C0hGpAcX7uZBlD4UbMj+LWU646R+lq82hT6M1CZW
mD8Th4bQNzrKq+uX5STLHPRcmhdVzThpCkFEyML5EeB3I0DoFwSoxaXYIeQYxhRCuMwhVaphKzL8
HW5poFHFmTaiVg4IkpsAMtHDvAKifCR0lmQP8sEPFyTfUvE71NbbraY8z/D5W6UqVkWfXd40P5k0
Za8Phwl8xWrmNRNmJyfQmQbfym1uPsTYBnq8efun8AuAb4DOB84O3p8QyQ+tH0+QvLMm9uEC0k2q
6yT7frDKrt3DOrjnfvtqg/Hqu2km98kHdqam736L8v4El0ArZbg/hDIA8o/f+buf2CsawTaXlWBF
S7hNpVuixlmQfrvlCj00FDfoQ6bvKmcA/yf5hDZL2zaErOythR0pnQWxxPsaUgsZeHh6L5KiM4w9
MKYrwAfamLo1TVYZE0peRJ+Z5db3r1zxXdEnD0bSge2Zi2WygidVv3O9Os9jvTqhnOSe0aqThAKh
1r1gawUQViauA2df32ZPzgMEkuBSE1XzII93GnFpv4wmuGgwQsDaf+QaoEuOZQOY/rwmFh5p1XUS
WZ3Xzlmrg5Bh9QGSuyigD1T7XYwPtfuIrrvAc1keixI2+5zwhGib9x+HX8va8ik/wenGq/hegKeL
M8J7FItyzHqfZ9yqaQKv8vEbNe7doAAAgOvF3uQHDW42NzMTioyON1lYk3c1qAuEfGYyqjxTXTR2
Pht3YDS6BNxPTmupOc1YJxW9OqBM9BPm33ErLLR1dvlhuzQNqvYCcPS9sWlwMDlRsiHXKzymXYJ/
k4fzcrZMZgSMmRRungmWgWUtx32iIG1i8LVHM3jx2ASv/acvcKP9/FyjRnEarS5QIDPkw4reTvKz
VCp2tfBocW9Llcx5YDJLoHeTfjuyC9cC19Vfa6LAYO9xTB2NjiONiI4OADTi+PfPBrON0RInI9HU
EFS2RAPgRmbip90PH5LbKkS1ItMu/cEk3918ofSGzz+ns2j3yQssjCjL1IxKjTsWgeUhUme6BcRj
WhQPE6diwuiQlUEXpWV6tWQSvTFqLVcJ6d7LngNyhxrCBgH6+HmXBbBQ/D06xsFBQNtvgPgAs31S
np1Og/cWNrgdgP8nVmFILy1wRq/AfaK/uwwq4AG243VwwijVCk34X+PeM1k68t31P+Ph2t08bN8J
RGBjvGufa7YfFFImIoDYiD88AhgZzRMd6JRuvChE64WdQ9BntssYo6//9UbwKVHdXrzQGcLUF6hF
cSrHI3gKERRvfq/1rIADHikvYUu0OwZE1mWfV4cdLw5zFiINYISuAE16RW9cp5YZ6RtJ3HyAWdJ6
SEoDRQ8DUuh4A9Nd8iSHF7qMXo9ISGYQG33gSPMD2RyEsy4rvhYpnTZGPObTa/4JRj26+P6Jd+ff
sQOfDGhIIsl8VGLzr3DYYGPY71cT7/DKWYCsgLoVuWPADkFWSuIQ+tGalsnBAARaLw5OEJas7Wyn
t7H89w59MjGYFGvgcc/upLj+Um3J1/dLu04sG/kQ2q2GiBNVjBFMR4hqt/9bAf/aqgKwYVrWX5VP
Rb7pcron17dmz+ZZjCdHFjh82XyBmE2mp0dnBlssd093WXlTchjCwZGCATMUh732nmSjWJ7HS7KM
xhumcX+nGr3j6fwc9iPmVvKZT26BkaytvIEG9IRjp/yM+eeA3JJJ6SUc0ZfNy5/KNiQeLXZE3d4K
z2hqc48PsZjeGbgD8l33O0m3SWiU/qVkIJJ5TQHihYCAxbNPz9Lo9zotKKhXet+MB2hkipGFT/w3
TKosQxJPU/OnKKsTRpe/Rw9k+BrAHAU0hbE5VBi6X9+0+CjGDnSnEYur1zac4nBb/tL0De0ai4Yy
C14Oc8ze1Dblt1VtB7TRd0vkkPjyzp8LcHiySPr5lsBKvlyAuObGbspY6hkXWztwsKqghmbEdRMO
u6SfWT1/Czg+PkvBjnNgKwnAgEVbU47B9hcbwaSuy1tQtaaZ8fjp+/EkmrcK4m5DqyrVjetLpty3
JjzkBtSa0wym8+0u9JANPm3SCYjiiXj91yTYQsW8nYKLk8FMbSvAY+4i1wOfI43izhqizbR2PO1L
jq2zlfonRy7kybyMerwXE2ZDodyK+puoaFoM4dCJRLZ/I+d2E8xmEUpFd01jnkxXOOs5jG59JZME
KGfwooZ2gAfVQKRwBGwpCZ/QtI4x7730noXLpGmZofEwe9au14Wi6l6a3FI9zjATWiBIs5bOh61L
aTiri0kXHFQZ7SMVoGG/DWc4f4gMOiyUJ6M0zXp2tMk+SNgKcGemG7pgXsInNAsOr00RXrgvheFO
xEwx8ny6gqa0nYGOygZ8vYMnCRkXAaEP/RfoRrxcTk/b/hoUN9VreFZOvOMJHYOfLaSqQQ4oLB/k
OiaivqawPdCP3esZvqCiFKbLx0gFn4qXgVeKJcJSTZcEU3EkF09O4vLtuHD6buRlF1GLClkQG4Uo
WVt9aAFLmDrg/JVfsUX3vvxBc8TGv+/3w5jxQdjK8MMgokSE/4aiAIzgX3VBIN4WlKg2PcsQ4FRh
zBmIWCsUHoURipm6+wIW61iuUZHMvNovybcMf5VUXHfKwkQMaQskxyWMKbr2TMZWMHmlrfsHTvHS
i0ZW82AaqrwuiSjkWOe4fLeKXd9jqgNWw/GEzjcNGuY976xn9s8EVMyY170uuKNz9rVN7aV0DphT
tSYe9YSi9ecdrdwr6int90ivISxgb/rmR14JrrOgBjWZxtR07zA7SoF3YB8zlEMTevm0Nw5ixeXZ
QJ5YqJBH5blRbwPCF/HjPOJl7iE40U7fLMDm2Epu2NwTZrFuVA5uAYzZ3Lb5NvYnktXWBm+RX8kM
Of52/NdhAC9tgWIBdXSJpZlPHHH+CjfCQNduOkZNIuGqTkqrRAO6+Fj+Z/wrDj4YKo8fY+G+Iu/G
a471SgCJt9ztfEfXNxxarVEtzXJiwkx7jCCeIDOyGoFunUD2Jkk86ezgXAnohZuxeOsLHysb3ryX
Ul8t/HTn8yfHutlSzwsVWEJuV29WdF1sS1P02qnfgxjdQ/U1vAy9hrIe2ADz2mZSbRouFqJF4Uz0
6TjkG3eIoLPgtOZcWds05tLcKkdnTH4zu+KZBjTnGdOgJ70WrSIOzUwwC/64QWmBtjQILgmJ4NLE
FGSMjiVNuruVDaLUltHyHNRDCInIF1pVepSoL7O8NgatuivYhwikDFrzPRCz3xpMB2gDvrfNZlkh
+gKfmvpI7LX6/6gur0mkrJ57lL7p4cG43AfPWMq3C2yed0pLLvE0z/NDNHll28QBlViTJG1e1Hzm
s09WpNhHz8ZunXwXVup5FO9KA5lc6LXv5yF22wpkF5RwZfMvssHKDrP8BTiutr8u/1LKSFprdqKh
2lAKFw+zgcCeeoti1ZkRpKs+mAS7pZ/JnP/XVa9UdLOLOMpXi2u04rzPujzkQLtB2Awqy5d2C7Yv
za096DJqq/G67EasVnqmoEmN6netfFaNjsVb8ld26UQK5CsVanhsEDiSNi7GRWtk2tsr1f2Ihq3b
1NmjBSY/Emo5HNxOCYZMO4CVkUFJeNcnKbpecfnYGqGgAIVX2KWIxGOV6JL+7GKqEZdR7o+cXcIX
4a1sG1pHePKcjoqRPPZgtY526F5ij2N5052meXCLNzIfMmDPnvVOaOYyvHYMRu50tvY+BDX4TRzn
knjMBUk1L44LxFwGETc+zYgjeGmMNwf0P5F34ue3/k4U2UyiSxRzdrY4XHMvhJPSTl2l7p2aOz9d
wN4XWOQgdx4qfqMKzNpHwyrLQAsR/jVw76WDhwLMpRctyX/l/V3syRtg4Hi1fvJeHWaLePs00BWB
q25k5lQIDn4VBgpN5PgY4xeF2dCBcGZLY8IPYibyY5xk82axC0RjQL2aVwoLb/HZr7Zj1Au8ZNAi
gHBjFkySxSpjhjt8KDnQ7lCjTcwCM249LuWmt1V3W1Ay9JcD65l0JqWv6GrbZ/PU6hVXGpdqm2+n
2Fp9dT9kxgl0BbH+QQiqlrhcx2Toiihcylup+7qXqcPRM00y9PDN8PKxr7oXUuXkdd5dKP7FvBSh
AxQa6z73VbtFCs9nQH7O7U6+xZpds0HT9ZAAPnwWz22+BfmAbcRp4lQCrsLJ4mCFlVmV8jCfdZPi
x0PgwYnSfUEZ0pgh4NrWjcwC2DUltJdb+SZoaC0jU1MaJOSHi6KBhgNRW1SWIH+PePtc7+h5VVoH
bFb2KVjZ+UB38/0zM2Uj3i1wuKl91mcNHjpXZcfV6sIeZRRAcha2SQNFJJvBx56x3jXD8VBGN/bU
UfW6gSGyKxQZIMT6m/3SVaVIYVKC8d89WlRFBTTgkFTgqYUvjQyciTs1EKITXyF6UQtbbR3l8+Wm
LXbmDLqVDUITQIQRVyP5eg04rOGA9SDKpdIf+4b30O6RxVGwoeDIo8vGrG7g89eMTmG6Cq8X33Yl
9Ur9nPGpW//01LCyNrTys4uk1uy69QmcecPqFQsXkwUCenPGK22tnD7q9QhtAKQxNie01S/v81UH
NDrgClAH8n0AX+fYbFahmojL+xSpLmE7Hoj5YodQisNg4o1B2XHNXVu2F5YOEV42g2iFQXkW8dPw
/W6QVgMRd+yq89azEJSwnKH/VbT1ri+cm9LXfXWo9rMhn2t/89hYo9a1xCfPbkkHZSCffqxj7Eo8
1NQdBs9N0qNvD+ds3kI6P1N0l4QucZVdG2B+4e3CJG4KYf2jRYwUIqajcpiO+ebJvMFDN1c1W/d4
JucIVxl+Gx5vEey68qjW9TjJvDS2FothFzff98XKfRY2DHc0vwOQtNXj8FRignO0fwGRaQ/NX2hM
DFcro+NIFX5Jnv3EcPWUaRx5SuSzWB2OeRvRwNlPY1kl9plIeavV5l818oYQ3U0MHeLRXHq+4X2R
WXkuUg0WxEBO4ls3bEzqUik7RTNJmd6BXmaoS0BNFjs2iImX3qSSB6mgXA/KpN3rYDLK1T1x8Hb4
BsVg1J2FpeZrw8ITmuwP6hMj731xaqPFXq45ec1/f/OHBgCOG7Ylmi0/Q2I8qLJxM1wL0RCUj21C
q56X/WUW3eugU81x5ZShcPvTTBnx8Ho/NWTmhNlhCJS39jU3XHJZDwDblbfHUuomhMSSjQ14azog
lQ3nhTjPma/9r98w3u7vsSjNpJXxzl/Xd6XozSvhCNT3zVz7Kqw9EUWBXMRThLgzfAAR9vNAGCvt
Y6PVQcg0L/jJMsbvSk9hzcuwS9hfcv5lZUMss887dWn7eHx2e2Dzu9cwgguALLcdU9heprYYxPGs
qavLE4YDSU/WnwezP/mV7zLAEqsUr2/IMOZetYROdR9IXt36iY+fYTUOhIZECL/rgHpDDDrH9F/w
ObdChgYSsoQzDKd8Otm7XVIVfj4l2VFixyVMeVVwYsqEJLFe7slPIT3CpVIEc6nOc8Fdw+b7+SsV
LB69LbVDs5h7vfUc/aVLtgTQw9Wdfq11LeKdQ9/tFeUUyuFsE+x58po7yIaCxBsdH5XuBVjj6xsx
o8ryG3I60QQCjCKZCXALfQ8XybK6VG+DUZgp4VKGiMKTybc0aoXB6OE72m2w8C4GdyRvLh8YZLfa
t2eOhVYcS1BPUypUizaLvSsSjjNtamk/EZV4bx27yZkfOBvVTzP749eFsFG75QX0RBUsgIyHqyqo
2kLHRPDNWfHPvXJuVOrLty0DvOpfamaWEYCmBv3iMny576vxHM5cjBNg6MdNzi5uzBU2kdx1XBsw
i28N3x41qC0K673nWWMD8A7S0Hu3D7ucTx0nmQ/+z6AhiUR/e9IBR28gjx2CMBJHOu/xgPTZI3QC
4xX6CPSdSp7XRNy0icMuablhbnhcic9stso/Z1sTT0HnZkxFPEsw7Fwk2cQa76LpshM5pYBnrRvo
1n+9e2D0/DQZIk3pZwyl8mRY9teLGBqLFbAYelwLHAVh8z6oH13aINbsWHu6lFSGbyIMVtcg0G3O
bEYizdeFjzZPENKGOCVVYIgW43+TK4aqMRFak+vRAqeofOMbCKSLQQhNCiWv+Jaak1FJ2SecwUc7
oQr115bjHc41i8jLgRfI4/2Zl82xGkx+7y1BuPHK8VNrFt3ga8Ma1QLCOEv41KKL1TpI0RcqoYrC
lVW/nnx+al6EQaRm/dd4C3KpYs5sagqsAKCaXa++FP104+kYg8BnTFIlVdRYmYNq+dQmJzpMM8E0
wvVLvmqulP4VD5mhA0MIhXJzAxUpYf0Ij/kBW0vee/dHJiHLqGs6Tr7C0Pib+iSR6EDJTYnUDjS0
r4tF4Io9C0LJR/w6zCry7daONqcd2psQVMMPpnDI2NpDxOSph1r9QMn/jnG7vfKF+hz1GVza2H9P
2jBBh+pkdkDgl0+SmvJSdlVisWOypWt3COA3dfN0OgYW0JRORT1deUKtXxxV2s4MLPphduvd9F1o
o0pgql8AIbj8EFOx9W9WwxkXQL0s3kkQ3tzpEbwIlHXPioQF8EYCu5QEIDrpACcESi1zQIARE9q5
dzyW5vsaYHL8dr5jgm1wyIGRZl2C9AwndSd0xeJsTx+oigg6Khh/cslW3KPYFEga4F6TCzNI45CS
8SWU1akNYlGWD40Jeez7EmVbyoLN0t7II1bdFTHsdEi1+jZJcDIM6Fkmww+k6eY/dt9xDcCzC/Gk
Tqckt0XuL6jeX3CQJA975sTYmOER7Y52r7CNxQNHymQ6QUnlOjYuC0FUoxW1ZvnKqVfiHDxrCRtr
We2Fdxr/rtJnpkthk6MilkYY6yYBqgo7YClVEIfsiBpx5PF+HwBEW8a4SL6Ezhf5nhmpwt3DYhKw
brz/H4UHfhLMbAIhmha99uQ1MZMhnYkPScEJAFneqC0ILvUuDOXJz1HQlcv4WJmloc54cZA4mwah
EbhBjSRto3CF7XfonekPv25xQFdJJmxSmxkQmBgAamtZS+OcSHAQg0vXsFV11BhoBe93cFSB6muZ
4r5iHyx059iw5hcOMJti/HZhn1qDQS3NmwGFPQ4GBOaB2ppxil4hjd/QURA0UXHtcOVBw/Prauvm
KiGfAMxQ15xS0H0LiZiYeAiJooxwMZAZ9Q6yuzfbU6rAyGnCQjsMXRNCCQF7WoDV+AJF9oETvC/z
q4Zs8Wgzazxifhjtk9zlSHjhkYcQCV05u59jJ0twfAp4EINdK1tuiqldxZtWBXysaBSd5NgCqC27
MoQOzqUcgs7B8h0SMeKS2kk+FJn12jKQui74j4Y6YJiGVoyXmzuivQ241bzkTkK7NCsIuhHZ3ZeL
KZroQHPEWRJqggEJiVm6yz48RjQ+WARKYN8pOds9PhtUUoy0z8QPoIb/lIYj+SK+PPhjHdutQ8lF
TAObIu5V12Tohp5iaFO+LkaCC5BWEgGqGsdvtVfPx7HaafvWzQO5NN6E9BoYQ6P29/QrvsRLMS6X
JLECt/w1E/M6v8fi/Tjz/mvfbLSFjRTxK9m2fZR62Lf2HneeWtXlCpDkN0n3l53sSeqaQWRsQVgr
SZMDx3fnPVnEISYcBbLZNeqbGdk0ycniq7nn3RyFyj/q0/wE3Q+rI0BJEcDBRw3UTBkiEPoiOuYl
W4tkhV6GS2YoHhu+u1O7D04iihnucwmB2iILjcg68cQ3tOjdYM1pVHERgIUNJdDPlTQyxkV21/oQ
m7FdSPcv5Jm22jNDDciReugVw7UmfnhWcoVlUvWRQe3OFUk9t8mpyr25G3V54ybPuuAAxK6xh10W
vsk3b6VgNr32zmcU80CrSW4qm0kJGuiwcWZZZO+a/x3TA486+GSzkCOxU6UYWoiwpC8SbchrpidI
p5b0fg6N6y+hUqZfQk2OnBURhyKG4aj4QpjLrqdR4ahDzPcQ7g9XRKs+LP2VYcMdjYrympZTIlNc
pL+UeIIcMk/C0+QsP39cScWCvwfcCNiW2C5m1gpC8kelviDdf79VeQpRU0bCWlj3OabbWlfcRGx9
ilXmdkPBnjCHZdcJVADdsokYaJwaOwEZaoo3Lb0IudsgnnxyOJsQIjkYBunYzI+eRGC72Nzwg647
TrDco7zOXOoWQjnIPChKAH0CG9HRap/9l3PYwGt7R8tEEClxLyHrrvwZ1ulyGeYEgYG/Xm7vVdUK
t/l3k6H456YzKCAXWyHr5V66OMVvxF9c1KZ4JNgQS3iIw9WkFr3DYRqfyiXtyuHe3+frblB5KavI
/8Ko7wYjcmIX+wvHBrXkPbWRPzLXNIvCdrxBNZxFwZnnnoffahmjvwW97bzRTqW3gWuXdBYLjI2E
FP2XPAjxWksTeASjg9PVfsXEZsf7UJeq2PyZsp4NLi1H2b3X2v5tbvZeim4WgH7GcWnTIEBO2XZD
YQes6x/+p5KODxgnXVi7UFSvaywk5crfRKpehFQ3bfspNR2ZpSXPV/X684N/sryFQblYcIdjZ8SF
I6KRifebBuIwb+MmrTMMsXC8HfS6jZ4gR8Q9TjzypGnyzMhKFptmtHADRBC+m+7hUA4TUArz/lyN
otsw0wFZldKKPGdxWhyg1KNtdHRNxDsAMisUa6ib6M3tQmPBZBRE5Rs2946ANBCZUjoWPVLqAzLO
pVXYBdih6i2R/AnefqsXgKy/NuPCA1pc7UJDF+Yg8q/P7h6+jtFcV3VKqn5rDwSrdxKOQvoHffZh
RJNofzWXk7iX1NBuox9OwZvC0Tct8HvdIZUK+H1Zj5WUqR12L+kSUza62VNbUs/6Cn0XeBL5ejsw
anh8PNfwoTWuAF2Xs8LUB6OD0QGjziCuwEbaJzYQwOGNvU+XUsmJ27WtZ3PCdL/AlDQnT74vOnb9
76xlTGU+twgIkZop3SsDDzWze5ZpbNHlI7sB6IaKFmngQsxSkwjqVWvmLlnZUv7hwfI8SNVV41n8
pDcT1zt/QExULqhie5DdEeuqf63ZuAGHzRx97sFnmfmIe3niPftyGykUq4judozuPW+QJ4egOCVZ
3UwlgE4zRpdxa7YZHndMe8frD1dugdvHckf6zkG/nV4uUDEg22e434sSzUMVz8CibJgS3EWnDxES
jE+sh8a9W0wHEg7E6uRHR+mj+IHE2e2405IoZhvIH1FknjFkmuXnZhhJ1Eee3GcevNwIwgPox17o
fazzRcPyVV3eAJgNgkrJp0CECc4GhUhFD4zUC2NeQULOWVSU2/mRI2RltI0PQJu2XbEXZBKzK1hm
ueS4KZYCccnv8mYZHVVnZtARGl2nXMtzeOjgBLo9clsCcJJoLPdSJ58i6aR95ccN9WtiKReRTTzu
qXtdj49ociV1MPaaCbBQBQ+KinxJgKdpOPVveIQHl5QOFVSBUGo4ZJcTlQ+QY0UNG8TnGF0bLlyB
ODRdr801p7wfMN/gVQj2JwDCZ8eZDkCPiQ+9eGy/ijhRrBml6eJ1mT87E+Hi3+srQVQxy0pdj/O8
3aNN874pPlzsW9RXKsx5iKjzXWwftwPv957DGrtQ0yF7QhCJlZNqIU8SGN4AY6BaY3M4GkEO0A2M
I8lK97mPv7ioStHEql71XWjOD/M+Y8eT3ppBLAMwF2ujfdCy0TH6Brhj1lyv4tNlgEEcfvVK2RNp
U45tJ9dYEPcMWR2g6V3k+7sAzp80Vfki2+fGz9HpZfohHLk3VEUXoYvgFZKLKLe0NYE0mAj5CShE
eRG6Tw2FhuNLoGIBLlqtpgtmELdoEbd3A/FctDSslE00zM4RM4BoqnguFBts7kbM509KuX/JmLo1
Q0TrtPP8o+9lbP2XXuJI6LhGZbEq5OPkylFJyVWbCLhLn52N+7UzAXmmlSjQyMtQGIqhuoskJGkk
OOe+cr85YGHQmg6IA+uqrIDxWnxlqgPktsumoKA0Wq4aff/IEK73FI0kOgezY0hLsW05ijYZ3dbj
Fmq63dm1AarmV/4uFE2gd2KXiZEq01IYVrrKM6C1rkAng4s70tJyF477r/whSArI95Fdk0a5QnAq
NQJgsK/oEei3ztz5BTJJqRliqsVjMe07qkV0BhQgU1X7k8hbMG+6qgy1uOTdV08V7oeEpDM19a8N
BhLu2MkLnaboCjSTiRlOr5gJlFrjaWrziypqPT21brvuBHmtj1vgifTW5XPfvpz/Q7UA8txzU2m3
reTZu6i94CBWw1+Uro+Byj6Benh85QEzEQeMX0c26xVxOOwiORCmEssreh4MD73lJugsCw0yrTYo
cMhrDXMZmxmSEj9aI1Feh/UoffumuMn0hxddJDNAQbsqiRvTaEQeW491wNSWJ01+Oh6ZmAnM7G9y
+aws9Mju5gqBLYKiEflBtAVPpMFkmx0t/KKVbCFGr0P65XgXHmePQSVG3FoXx58VZgIU6mC1vI62
vT47SlmCYiGnl+vScfFSACKru14f3e9WDEt8zGxrFWkA7RF6OoiyHXJxq51dxSrDPch2BOvcmFJ8
YRq75GmHLBMs2nL12yhIMzfXycaB3AkYntKSabKDJe/hl2UAtaMCJ2p7kp8yCvigxv4xTJpunOIb
EcFDbpeNekbdq9ZGlwBQbCMjnCRIxWjpTp/TdK9ShJKmc78274QUzYFdkf2yjHKEIkfoHFkUO5WJ
bFMR2CJGxCea0XChHh+Dhke1Wt4EY1V7RYmmmSEEZp+/Jh2sY8/iD4EIgQM/EUw4eAiZTaTnaFSn
8sn6Nv7YEeHc9nZbwJ2TeDYj124i6jMz/F2hcotVOXM+BqSdsLhDo2I9mlgOYNfy6+slelSDY+Eg
McOLxOHogw6bq0OtAzBa3oN6UyytnNB2Uf7Cm/xiHTETJH+ZuDRXcsDdgZK4mWNVAaXiWVqX821g
swK+U76BMuBLcf6h4c4f/KYSHD8j5lrOURlVDmSwyJjV7s2qHvTP4Qr2WYUESvJCkma0HhI4b3pH
qb+iElMLUmxIsD9TE7cBICUpDyF0PrRJX7TfrO5nyMqYycJSaJxCdUsxLqha9Sni8aTN23VVGO+h
HuxNxvr/YSUV0cMcj3AhER4PRzGcMW6QYalZU4bvk/O9brhnOf2eAYg2vmvNGAuLMy4IlrHDetIy
nWQEL8EfO9Zx1Nz4aoDDL6uwhUycSqscroLULgoyFynvwoOmmWA647gxbrUxISQEEQ5HXlimyQxj
dM+tMq5aLwPb33s1tPjOz5FoNKygp7Arf8eB96BcC2/Wii3heM7FRphNQ1YpqMdhL9TrBT60IFyQ
EocHRLO5Oru/FsDQENq61qTOFZ94TDepl8XWeCpM1olS1OjRemAbu6CYMnQs5C1anz3qgskrC0Gy
MEpQzxbQetyCeCZwVv4QM1+fFBl7IC4YJL3ZJ2LlCNK4YE39gOLaR4DsRadqYX37VTSm+z6nqtSP
fIfz5ACHUXj33RRc8zCSx02i4a+YlIPbRo0+p10AvDFrWHGO7N4MMcYJMv/mxO5M8xUXvcqIp9ls
TMmuJ7l4OhzQePtBkuSJjCVDaoqU3tdXWmlyPJOs4VxPxlY4JLqiTWpY8dSizmyjSLr7hsEmiBTA
ujHGsEDDqlZ3W9Lc/ObWtyuSAdS3kFNO5Lql4tfrZGKD+6K98kPAZwkzxS1ggNbFjA6T2ufeBlqh
FX2b1t0br21JDS6Nb49L+c4kerO8JORPdGXuv8J5aDebZ5ohlhiQHUarNPPad2hFAjH0qogIhIzi
ZXtiYWwco+66JL775+mI/5jjYsqkOuxfPoChaA79xSrOCvMLNaKYDuv1zoApCDigWsPLcWUPEOfy
JsLjwhaaXJ+gr2v0jMaWY3LOpWpEMqeGHsNnoF6KaRVVewwRTOHpK6q/6aEttyh7Sg81HIBpeCu1
kkn2nq1y9oYE/mfYzsedUYimQaflx7KaoXIVQZrta5LUlDSTN9/fWBMUB8jfXMq7onCBGHxf2NEf
ViYD6ROCxphWam5ZapsTaLg+mkKGxvYqYi29/8FbMgirBKfTDL8OPBVICsImZcdLZwuSS5+x/Lin
oI/KYyLHdcgBg21Nfpz8oZBGop9gJU9L0XQl+WyiVFOdZa3kwj+2t4GwVYnuqW0BmU2YdTxVFSun
dOOKvulIiodfWDg+gRDmydZjsAc+oOYV6KRyFH6xviFa3GhtXJdw/KaXqkRbjuqzMS0kuew+2fgy
vxbtkG7fXge0VM3F9f8MIn6zlvaaOqXvRQgfQdtyer06cjLtWC2SbQ9/x9q6goZ0/bsc2m4pSuE8
I/CsfebdsqCbF051p69hDxef63hhsFLiS09OY+4PZ9YbmLz/77xiaBT+HTJvb6ztzRHh42xGpCr7
+OopWvHdVb6MsragoCG46lF4EwdaR52B3RXGpZa3E3wp9A3HO8dVsG4kdQ9hS1oJvIc7ZtLyBzBa
ic0iX7VxhAt85NAGp2otPpEUDeCRPjF5PV5MiJZGB/W1YyAJUGZ9s/7Hmvsa3nstdaTauCDNApqD
2Wj6WKnDul/vTuB1e4IMvuUzENAXRG+7F0Zda4PMXKSI/XA0hL4iPefB6Hd2+6uzr9/bWM+IxG6Q
hgeJDhoFXoKmxcraVMNSA/bcATgwILnrqmVb7NzUAWoUbcVXd9jWaB/b9aRz8Fp/ei/676elEzrD
iRY0h6X3zWLrPu7jyCiXzXvIu3/Q52ZzCTO39pI/FGQaTJgyyhrdOxnVfHQH3qxCRTPByr5Uq3YQ
CZXAkIa3pcyaOro7lcreRbBzgiPCHsaIadGRhXU99vd3Vb23736t+gA9BfIOGi2wTGLTNy2m5HqS
SfIV/nMPC4PpKYWJ/01rn8oDJSfT5ojyCMk4HT6sd0GsRf+gIBcjTNKvXiHb+jRgik4CNNQpCGWz
0Y8RaMD2ZiOSKOdfk8tVezIn52QiVR7pmD7dgbEvyHjYchBiRxAKAfD2oWQwyQAHOWObeKdKB/8b
hmD2byxnFfJihTt9EY8iqFS3m/jEeV8B/Qk/CwYJYBowjX33Qy0BSuzwKrlm1u4NOk9ROqNdy33f
Gx2d/P1QCnqgfCa0n8SsSd7mIhI99NsGwrk6hLjqHfnNv5zIECS29iEa3sYbm3ceHscCCjwN0P0y
KFNsOYfEMewXfRUvW9kaQHu7BNBVDV4G1TglBFitGesgnq+M4dq4IyLPTilKIaJukGQRR4ARwfsP
CzM3IpZBFZwT1bYrXCbb/6lVh3rQAnE2A343tqc3NvjmCUQdJ9h4IazKDRvLuvw7+yvTCPqQ7riJ
sKeSH9s9JvijPFJetiuE4u+SMRHxlFYhaLjGFCv6ZyScwbGdXHnEtzzPKTXZiQ5DpkdsqLlRU2Cu
j1QbUsfeJsu3pvAwkORnAU7MiPw6Xa/q7sgQmZRZAq5DIb64GVI4p0ieuGU1hLV1bVpX9ItPS//x
O+fXBHcBK3RCmMcM6OVJNvgAJ/1vG7m4wyNP1IBRmaYw3/K1/mOwll1cH4kiHMPLfeLkr7HL55pA
Ai9dqbfHelASLi26o7Zk5HeOMyiQAuqyrK2Mr/DHjpBVh8PXAZD97VRmbiMoxan5UosC0xgwBCKo
T/hPTx8Q7RiYe8coh6fEtZHtyf/W7YWDxYsmtEnk5ljvNDRvFdDw84+yVtd1kKPo7aK5mUfpy1BK
brUBe+sb+04SbfhLRZeSRBvDt/rRYFEp3eugYRFf4jpaIqjJyxtEzkqc8e8yvB8XtIE9rie5ormr
G1ZChf8qMdz6RP/w3V8Q7sLy9KWBkKvwaxWnBQnDKfef7fybPx5djSOwNt0b2QDLVNGY0QzkWH8G
BUZla7/YRPInzg8Qh535JX0jbC7xOZyZ0yZHHE7PpNCDEf74H4zSaStTNrsX14vzboukkmQa4ws8
78c2nBeJz43sEGcl6N0cGanPxmqPm+5FdIBTdcgaAwuJG6mg3WTKAe+tp/fd8kerlkB28XaC4/qv
r4fBs8xamOgvGEV9olltQdVllXCwuj+w1Q2Bl19J3Z2oFFZuJ2IJoGac+aojRN2sd4si6vPKvH9q
oOZ2KQd7UxGob+AMoHTbbSNm3zUV6QpB60Hbz2JxGyTwQ7bNUygCuQFjgtrxeDXkjDZk/HeX4pTI
7jAZGkiozKpVZSW/+pWeaBgAUuk6Q4uCcTDfNuDCd8yQLz7EhQal/LScyY8+p3mDhUyLrQsSPMoh
+EieriJ8sWB4jKxy+FgYB5mVZrFLiNVsizJGywqJvgGGllXFW0PS1rzRAONWVhddfZRSUXpp12HN
bWtfrYuX9k3dTfiTUI+IKjC9Bw6SpZfw8uiQHwQ6qfnw3Dq5TlkK3wekD+poIJzRao8ab0C/lBq3
ajq7SeF7PogzFB8PGAY7xy+Z8igkPWGtlQGhjf0ZL9wwnvEuScNCqTLIMdRqMTbCHylre6qgwnK7
SveL9gxT5Igfwg5kTvQHiGcPKEVXFDkhaQd5DtnOLZncZ2TvX7qSTX9Q68zj7ZIs2GiM8OP6kkIT
/qGTozijFXha732GXV/gddf1vXPa3NDW5i+AqUIGy4nrB+s5HEE7mvC0bufdKZLBTwYd8sP6zRAN
g0KxtgVvEQSrLm3PtVFXR4TlEjSqAOUCyvX6d7GHQvga7V4tAARuO/7mhXAfrHFRTnHYj87MNH3L
MLOqkR1qdIZbhFEyFdUzqaBQK4TdO61xzddQPw8IraBw3KPw1gv45jWDgInqulhOwDywGjOCmEla
FsybrgydinZgkU2ckFe9gWwypmosQ3SHOE913tNVheZtnvdKURStR1MSS5BpP0/UKC1UZuyWSCX7
ItyK0a17inT02xEXihakbtKTC/tEXFMteOVBjlPjrIVWmwKJhrQXsKnNWFyGC+OsUxb4J6eX8uXM
tAHE4ugDlVWXoNW22fxb2fY6jIralIZvH2uAWQgxMSKeWvzFGE1InXUliKRhN4g9KkHDG6QBkykX
LzYJQ26/XJGiQWq7lbcJKsWds642dVhlHOqZiFPAW5VXBdSut7TaDUwKzSswCecaRIPSNiVbHtaW
T3eJ1uyFs7QEbuFIYJd5P8l6E7nrLhAkPSOh+NeO7cxEvWaWLTzpz35Xc0S3bq9eiSSVjY6nCBrk
RhnQz0w+JqZbPyZYSipCLJadrHTRvPykNQDgoMQVZNADeZ4Mv8XjJ1zbAxqWz9/Fzg+Idjx+EWF1
UCONkeHuETK4VvXs8Z+fbzOG2Mq8M0aH7FJIq/Mog29ljTO5VxSXzq1bDQBtDYjBwkXynYLlTSkD
lFZDUDYjax1X+yyaPNTwcVgSQJsW5nv7x9qj25dW/PwA0q+J5Jv059UNtGMsL0S4zdGlmijfppUd
EF5XKL1GKrDjZseyUwOC+VYY+IyqerG5DhBWY/17MgdXh+W9cEemoi7hhm911Bu8mYtl0WQqky74
0ZuAIa8l0CbwGtz9CN8/Fc1PIe0DkKNt8U7CEgBJMuA0vD4Ct8kIDUng527cmLgHjszaBb5LV1ZZ
Nvsh9abM8RPB4SvuNlqvB/Kei4/mijzz4pX4vRMgEWPIuiFd0zp+dMhkie9Wa3CaKn4IhUg0bx1d
Gx3tKrTuE/34l6+h8pHZiTPSCpM7DvDZTwUIRUv22UR4XS/YQQwIa1t6IprdCsoUsC0gKl3NWwoK
dE4TUa6HxfMdUU+bLQwWUXtxPc573oRW+flTEWZaAV4+JGeWE6qpDp2l8XONxPAPt7d6Li965Sjt
l2MT9PafNTCCVGjylL9PPa9Rc0kA2ltsmc6K5R365bzDHkqFH3VdzSgFgDtq6eyQ6PIW0pXAaFka
jAiXkNCsIi3LvTLUQU6LXisD8zWKflE/BF3zI+z9GENs7d47ZZW/C8Kinm6Mf5qbRDJ+j3v1eWfy
+7bL0kObUoq4u4xd06pU2aeK21RHI7iDILsAdt1zObdxXs/xbzWZw0cUzrvFfKTF16b8WO6ZVPQi
ljiko3agqUJAUilaSwsV0HTyOmWRKsNV/wdqYmYOqJMiBefEgS3la/J1EJfd1oKtd840jvai9hym
6LqNd8B/FUUPWTXtWPMEATeUDNwMU+kCc6FzXxpsZaXZgc1ZTT/pM8bK1ayJ6ogrdxnijjLB2aab
2w3XOAyzcWGoyOQDBf61eN7Wq+I+/neFmUhESVgQhLvs9ATXzUPCKDMVcOW+77p41hAZs/mSHnj0
sKgaEaLcCBKGVepjgH/Gpcrd9OPN5dorMI+G1QUNDTZC/MuNuJJoqDnh1FKzDXYHjU4AG0GXVqzL
QizGyJB1F4q3jkiNYdOpYYPJfEHXRj84GozGyv8QhRI9SGWZTLmCKpIv/zSCtcxwt1bA7xksXpOC
iJFKPxm9QqTd+4gdOcO3DiNs08uJdz4FtrCCfy4TfOSZi/WQmJhfBaigSs8rEzjYgehfpT5mtgfC
mBtem3F7LIq7mYx6RJna4y6lbxrGjj4cbsr4bffb2cRCYEyicjfI/DjJymlX3QQt0LkHFiLLZUZ8
SGNgAE3M6IUIbd1dPA/yvksv5bM4yKhgviQQiXnXJW/ycSpDLrJtdiApOIrVoehGgmme9JwvKwY5
ySOng9yRnkMq2SSy+UtU6dRqOtKyzLuP54g55NwaQ4v3Gcri78WFxX9yY271y7w9mWCosKmQnQXg
rJrmYKvAkYOzqYk2Oj1eeb0fxGoripSxJ4izF/c6qF0G0JnUKuRXPXjHYfGsuTaXW+UQjgIgOYmr
xhRcKwfP8SutSMS4I+kWzd1Tt5zdnD9rhec9qL6cBnCYd7ZCCCM3evVCZtcuakEZVPpR24LQ9L6p
lYTRIzVfNEfUXxNOHxPAHnNBG7NdOz55TK1forbT88bdUkRedKWoui0TxjTgiJhbQkSS4GA/A49l
sxn3glfHaSPdLiNS7qAxIw8wMtV8wC1ZVgBRvdA9VV01/u/BK7aY59PqQIH4BfFPeflLcqdvveJ8
LMMUU1H13DIjOvVpKwE+UAQAThewStZCAiUh2EoZMS6M+7SyyhgwvUcJBFTsyOtnqUs2k2NfXSPf
OR7ze8BK07pp65ibW40npvkCgK3pUrI+7ht2HkcIMYmqGrmL12EJ/Mlq6s9nzZBPWWYn83QIE5ZM
7DgCGbC6XQ920SUplsFz7fk2YHzP4gZG827uZyhykvmeO0QgX4Li11A/l/8M/O98n63V7q5i9tSl
C0JXe77GO0cHQUG81XtJKAsqVzCvqA7MVBGJUYxVTntHODy/QEF1qxR/25OaKuGRo137CTcRmjvR
6bziFU79ZA+2GSGIohwm8bHK8DTeaGv9RX1/zVRL2xn6e5EUqqtcwQjcxU3HAXKW5QZBC0oPJDkv
THi2OY12n6vm0F6fX6vnRsI6SOHas98jSYPWngs/cc/LVKhRTuM1ZkrWjEvfeb/6l5CgfYRQD1AD
WshjxXlqL6tlfnzRn4EIk+uDJB4L+qYMvs6A6tXt24iO+yMF3dOxR0hexlokT33S0aiQseECsBPH
5PWZB2aQsUOTGNAQHOUZZX0LP2x5O1Cc9CyYHiYRbpkSDTKypAsrznq3gBNk3SIQr1D8en3C9yDW
6KcQNmWYarQe72vphaWa3Z2gthrr3/uTTg0fkt5nEXoNlwH5pf4LUqNt04r2OhRuGjVp6z0UKKqW
DDlpjJ3n1U4pWugVMD5Ya8d6NXLiOKCyEhpOgN+AP3gSMCL4+Rf3eh5O2Lepfl2vaSysiNAq5iKS
DE1fJED5kVlZJ6kchlF5kT1jzXzUhLNuEKhiMERD0/nYNohDJ9a+cFd1FMUX4QIt0+dax81imnQs
P0QEVdrk9lRgqiRlkX7mWdp3Vh1UDEflx5X8RoD4VUAwGGK8DOylNN7VEj3Na6aEt3jXJeP70dgM
+65zyIxa5x700SmJrkdx1Q5Ddm+VeI2s2qj/X7bPMrKphoS7Ob1liWc7DOT5omBCvRyW39F36llF
aD5rT5l6YirPmrrfAUsr1HGEQsMMiVVtPHZuKhmVH9yMOBFdT7bvS7QSVfTUAxanSmQGhNszxU4w
xn7q9MO3ESJThYbeexFi2boklSCWnY8tqaCdtzLdrSWy/Rhi5qsJI1FSwFfnbbIzp6MCSx6K7O+S
WoYur4Q0H0/B9c+B/7qG8Bhw7MUzurgwpbaVNMOinKfr8SpG2KicBVWapcFe0wHuGPvjrXvXyDeA
oo5TKvfKklY8Jis9E+pp9C3S0c91IB6zokPZKT5+oyDx/qyARDM2B8VBglSi8xagHPibpZ6/6P/5
+DpA2WcdJcQy77QfQhC6HMzzKcDHe00n30Cqb8N8nrinwZH0bLsUXiJdV7R+cFIGNR3ZGn4xtMuh
gccPaUiiKcy3xEoFDV8QdqFw/7VUlEqfoA5XWNqHJJg2JhodUTmnRcApp7niWuWm8U/orhyYgTjP
hCDzWs3f6kNLScKAKFxx/Uv+eAeq+xfBd+UHMVH6mpK99nTd2jsqznXdHxUpbYOvssp6h8w4SRio
K4qR6hCkzTNJ6H7REPFaCBleLrFze0Jo8wYsFXFGwLkk2OME1TsIiyrYRbqqUsBAcknsZIfAr3pG
fsY9pcRC+/dRFnWB5gGD6XSOmenRa1hzHLKQ6/nm+Vr53itN4EXU1aNXj0bl/gjX2Lts+12jvHGO
t7hBZ9DQw2ocxUH5PfEYWhJMvMW2WpW6F4fDIqfBjHbzHH3To3jl+Kc+K/Y11vUHSdu0ormKl640
/tVmdby1EqPPFD0bDFJp3SX+QqRaigBkl/Xz4D5sACoV7HJYH48svx0d4GWVxxi129+RvCHZdUgs
TMLkm95+ELvBfmolNeVRDzYV3j9ydR1zfIBrvFbbS8zQdoS0ytS243iPwaM6pjqBXozUJ4AUEN4g
/jRZMtBXLE/20GmLS4RYiEEtetCOqmT6eexqRi9wgW13yGe+CZZ8x5PnEOUNR2tYbG9N8Ps6UYTE
S0jFdkZkhU7KiM4K+NuqTCbvkGCqXnlpugVqkWxpcGzjA2aAHe/AZcBKiDtg7SbFLEiaKINtNR+Q
vB0YLty27u/JDqe+cvSkHVJSM4XsyObJKrbrDwZxQkpmRUWZ+UMo257L7LvkDMzcjvFYNrxaJIqX
rrnoNSwc0OcdvK6v+HrRpqpT499mFfof+y6+sfydYsOo33z/6J24x9iK6mktqyLoCdNvbIie8Kx3
DPlqiuvJBAZDdSrM044NKndFZw3oYHpWdovDWp7arJwxHLLFyR8zDgHR8+4DKWEEjxpjsFdp/SWH
c9/4rmIJiih45+hQnXnVw1h8Mh39fNzFANOq0xxHjynle3rU28djIB9ymylJgHQM+gcBiRaFJl8c
6Hu5HiGPsqWnxFSaZGinQGaWS7TElC+oVuG7Mznagyfy5GEyxQ1q8gcVbPaTV5GJDph/o3zpJGuR
JSwoSq75sPnWo/mTH2qJ9lNnvAnhqFZIWDEZFVbSgV2GDILgJe8oRX8afwbaL5HREfLBI1w6tKQj
NCjcI5l0EvPGpdAN/mssfZkDFshM+/I2JxvdW/QQd4ikJyUjPKhRJ7Byew1XNCdsrQOFS4SIGNZW
MkUBurRSOt/cuu1HCiKsM1zp233JSWxbGmk1BugGv2gmtC0IvrPs9Vom7pevRy/VZNexF8Cr5QMS
M7q1kOPFvD4uDOOyVbFug6PmC1CFNTZbce5bynr2lYBZ5kukG76uJtWfIaPRTvQGf8+BjVtDKnmE
IOfjdjiTduP0d+DubYDpXhCaw0Ry1qBJe482nzubeIvAW/NduPLg72mpLyWl33PhrJ1ErgkWvA6K
d3GL7ncRr7LWpluMfWVrTVWnR75943SUV3DaWB1M4HvaQde8evBeYHRVb6UKErNkp1PQcoaOO8Wn
B6aC4KkGt6mgOOnghU4KyzMtet/fp783HZFpbsouFYt5EEbG9mc6re7Efh8JBOmLCXgvq/X/ocZx
WizpsyNWqOSvkm0iP59do3gTKSOxYLdr4RylHkRiKdzfDBkG6rXHHgIVCejT3LpdB/bZGeNc2xME
zM7YArwr5qGw+EOO5+91uPP7MsQQcvo29CdnQs9rAi/pMnyfP7gftwtiHl+DzKJPATdUju5dgt1J
6rvHz+MsYfp7ajtaZSdpM+a3EFjHuAiXR2VSGqu4oZt6sdZm3A4K+r67doYCe4ULBNXDYS5bTYDC
V5Vq0IKkUNPLK1UGldb+ULj0BDqJUPqThGE1+xnmjgtKrOe4nh7iCsa/HhkcWLBDVSfBanm/WM3Z
bRRpLvCQ3K4v8O9gZcAj5FZZncmjYa+us+Z0ifow+EW+1laanrr0noy/VPlEdw7aR/4qNahfDpzK
Moh5Y7kWj/UzLR7UTLbGi3Qf1YudVT4Tup0W0ynyEB26S1g89yqn6qDW2UzLRP5LRIZO1PEN01OR
eSzsK8nELybEy0HpMNWqw5d8xLtjaxhL58U4XHUSBRgDtqULlgf7W0eyxlWrj+e4/aKHaMRWjAGB
oLMNr8IUSexyZKHiztmtk6ljHqiOL5tCxIcVDb7CJWCSUBxl0Kus7dVhBAQBBFPn3Rav6gVl1xEW
LrufUkiTh9j6CnnyWA9qMvRPQm2X7CllGhNEFWpKfoOrZOQjBcNeIuT67cAg7Am3w1GxplAML2rC
na3kgG3jNKZOVqhJXMIslQfaebH2natbNpyGoHc2RkluGTEt12lFehrE5Bk2mj7Nttwo/thdaw0q
j96TXYK5UHHvta+IqRs22FuIeZKsgBCiq3y+6NHFknCxIK/dSjc2kLHGykNcKF90fveUTMeiQWmI
V1t9Gw0LCX0h9H43RXcap958JcZgm3jZFb7ibHol7INpfsJQSr2f2XK+hSvB8hsaIx8x3eVWy43x
FjBKGYQY6qYMdZx5mS+RciYOp9oGxhQ1HJ0GBhRJkG3ItPO9NXcsSt4P/Z+wRABsY8ghcGEIR4Zm
VGsUyT6njJXn3tLIgwYkE4fb/B2XHlp41jGkIkLVgizhuRxchywWGXkwpmp42KC+HK9TtJKMhVpl
nSaaM7aW8PrTqhqi+CkZJng6DFJWU2dkGnyTaiheFd5hb6jQV0/ROYB0cgqWh7Pm9wSfSrdEZcsX
0eHAFAmy/PCGymH76AcoETAXL7CSjdd2wvfEgRauePQQe1+480KiS0IO0eC2D3HmpR2zCqsMN6S2
IYTfKDk90HD1YtpTEj9J5caFoDWOQ8x8BezJwVB461mfcNUKHwJggvGh9CfgNoBmclMj5KusxN4B
O2e3Cop89cRioxyWq7xBEMCf/9zLIRStw5cLR2MgblPhj1b/qsYqze9qSSF97uaun3zDCaZrBA2q
wPwrhGfM/VHgOTh4JJlNxrK4So+6PPdnZaDAbweGn88vgAar7cP11X3pAn/PY6aiZ4YL8fD3bvTj
52wZsW1jyq6VhF12pVDcoCpBJ8QJjgG9Br7l6RIh/bcGqI4vYbURP/f2KTTMamVpJIuDVauSaLPu
bwROqGYUNwCJ25JIHIx1rtIsLsLI6BzJGV7JbOsSxtJTH0ytDb9w10EkhJFuFaJscqSeSpYr06eD
8KVan8RBHHBeLcSP5tmtOClsNzSZYmfLBJOCArSresQ92qipNC7aa21afO0ugn5dvm6gZ39YEuMM
oS/u32azD3o1nc0BdigzaLujCU0vLAHNUlxNyd4A5aA+YegwtdF52YY7jFK3L6K/9FUJ82TD2M3r
B3BTVf2eEBcdaRN7WmByWHJ1Mf8zHhF3kgwmk0SfJfEULwy/q6QWYcx4QqUFXjaq9f7RRSMMgXVw
NVcQ0y1WaIDHAtULj1pmLUlSMMHTSb8Jes5lHM4U5NSL2S8mUQZRaG2euT96dwlEh1dSM6UFx+KX
ALq4O/ChXSQAnUmQQ474SpZgmwern1nd1gViUyGtwWEsSsK2FuP3x2DKjeIo9D7+sVY6+Q7/h0Gi
K6ConLNcAW4X35kroclt0fPkLhDgBhXD0FLy6uvNiEWLd/n6lrsnOPtTQfCHsGRNlFJbmxDKjb4V
DDeCe2RNIpBg7CvUZDjo2P1k4L4LaXc0q8FxAuAkiAhE7ySkbsjPtg/k/CwtqlbY8gFqLkUDvKE2
F8DhYBdksWT6Dt3YX4pXFAzqDjlaZgfM8bL8XU71M9LrFyYseEL2jedd7HuF+nRKKsQhGyd3EQxl
mjvr/iYkKq4yuBXXPfRZLQA3lMbLhYfW1NKZFLA99SbJvPSqgpaxgW/Ra1t/ThcVmkEttMc4lrNd
WknuK3NPgUurdN+NbptdZpH/7GPti02NtijK1mfWAwU0ahGVt26W/V5yH5qLjqBLXVuXFqPeLK7d
eWAyUR7o43gvQ9BfmW6Y/919nTVQP2wapRjO4rZmhhZbg3skLnss8fA7oqKykK7CS0c9mbew1eC7
OAeLQvW3fUntthP+Ut575kIhZqTOEK3M3lpCjax9OQl6okmEMfiGBmbCmhwoI5XK41IUCGZUDlQ6
KufLwAyRoWbjB6v17Gud7zxxIbCsjklXYccELFjWHZf8fz1HVXwGqbaxrTCpV5e+xV3oFkxtOzLL
CimfUYwwPfPZO5ctBrRMhYjMxFjcJ6iK3IsreD6L4s9KjMFXnIE18XlaOkSopqVonQzB3hIRdk3S
yl3gfJ0nZW29a7zserZ80fjP9EP+JbKDAlvkZENgB8gN6H0gzMWB1yWKtgBODoNTTd4jdahzhWUr
QgJmV+UONnX5o0wpoLNe8WE1Dti/BFMdn+hMP+clCqdkX4TUWT1Tc3LYt3vFVrJeuHhZ49dXvEuW
lulm7k2++QuBqsXsPwyPtIYgwPj0HD/NG2xzXT+OXtrhOt8usjmRUAlZK/8qBM/6anFMjVhsGeZn
IUorjMaRxcM3jR7W7WLU6Usrb660rsAoPvvVFFHZJHezDppJ9SXdhQhMMWIUFdRfJnH+aAdsd0Ez
w1+EisYHqDLYQTm35URWSVjTUoPh2Q0+79asUKrLb6YRC9c+vJqjqWKn378upf69nLxkOK+TZU/F
7IYpc64EiN0AXrAb+5DNy9g7emhVDC5VDcHCgFupKaQo6H5atxEvU0LZDTVlWUn+1wdsxvGOPKlc
1G9Zc1HF+H8KN3f8ALBC40OMTvJ9aVpd/laSkFrffqmftZyGPyW9NFdOE4DSPSx8VcPoilyiSrDq
1AX/3s/1mEZNiCgVeCyZxnGDfiI0YObPl0NixrG26JNnbuhvWRsirwW4UZCuNriF5g2yMZ1elnuN
mHnwZWal1pvVCcTHMeezvcFifPUuSHY6y9wK9VkkFV+YpE2m7orazriAXxrUJHex58+kfMvd81uV
gf35RyaidBmEmXChCkK8rKO3pXumWO9EIY+si2uxC+XJx+qQ45cfI/lQkM4OY7s7XvE/OD8IfMGn
WHf4UFd8zRJeqd5tL9y+Z1++GcRSGGHFIBMMTynGbnf6lrNfg4nqdxx1/uBTyc5sYWZdj/rdEWUP
NqaeqPfoxetwBpDcvkXeXj8f+0YsO4hZeyPwylcK7SsTuqbe6ExFQ+QVqALMj1G/aDZUbw5bOPZd
GlhaD7cyQatBouvRSyYvK7kJGvv2qxSpSVUkXKkz01Z2Qq96mX8IGRuKjubi500RZysTQGXxD96A
UDiqFnnxXn1eVQxgCegaYGZwDvyMFLrRq3uzXISS33kVabXEw3UYLMKL6LBXeIxTwh/oTqdjVhJe
zYExYL5syS6Zo3/QtWU2r+Gfe80R9aG7m1dCc9C5IfqOBeTBtpkAY0WLACKlcgRUrrsy1SDbKmNH
4T6P3pEaF4VgxAsfQ0+bsR6T6KJyJnDrve5iYi469V8hYaj6bZkuRDT4ZZLi+WVtZTpTI6T2vICX
nRmdQFwLiQ4EyygKoQd1BnUHBw+iLUJDHjVuyZ0ShKVTpc7j79/TFOiiwKLBKw3U6M9Zruo/wiP8
XLUwigdTNiD9hr34fpnjhaqUyNw1dlwNmAWO8tgLvrWFsM+qiFLtgeD3+16e9YAThgv7yIkt1XLB
p9b0DB1LXIAmTuh5oXo7K5dMNfDjbSHJEgu2Xocan60aHMfuZ2orjXMGWrh6xyV2nPv7sbq1KpkE
GfZc25ZAnCzYA16ej24tqkz2ykLiubZ1XMEHET1+CVtWKDghoo1G3deMtorxOwOJkwSj2gHXEFJv
PlAPTiEtCd284tKy0B9QWp3fjdeoiFTE1jV5wn4xFpd033r4Zo6N4YXsjWPI8ceoP9kHEKRciCMN
bOkrTLGmWy/BKjJXaZOeQiD7zLhRdUDaKzipIr3id7+7Nk0F1T6vwC/iowyJHg9JSoA4r8kDURmw
Pbbp/pZweR/mfUn09YiX7kD5jEehdzQFTtHN2tBF2/8t0+DNV7KChAMAYu6z9f3rHrWppUoQ6Jxv
40lbBFORKLcIu4xOX5sv1MiBVjLV6sqD8ehB8JBYCkFIn9ypzotuOXxtPs9JNpkkBhBeuV1TcDO8
O0P/drsHycyH0VsI7RYemHkfWkdZa6Y76Q2yaxN+SvkvMNdFSnnu1aUnCx3Dk72U+6c29xTzGefQ
cV79qRK1lmC+k5x9RUvcHGBphTvLRH4IOY+hSYqa9XXn50qItopmZvB5WvLBg7sRhYESqym7+t6N
wqCXhtFrCOOObnMsGDZM2inwBNfK/AIRwih/jusQ+9CWs5GR09TFZmDxh33ATFXQfXTShYsy6Iyw
JkikSgX/+MJD+3/B9W4ljJMRzYOVamtiEbm0NiijcfMok0rr8u/YudNa3w7rxpNnKTJLNQHY5MDZ
qhZhS+x6b7814ZCMwgjXB5mkB+mrkzh1CB98+8Wi7oBHzh0aX9VhoQvd3wKDMhgOL8G0qMNxa4Zg
ZeIeNDANSohexgrV+92Id6++4BMLbLYAzOy25ouLpd0Ym3RLHYWrM+HQ7DmVQgYDGUFVwlX/2cqs
HW1qSeQF7hK9NG34E59FjejdCdBzT/5lPciP9s+lMhJKgee+iHg13gb510AWxPI8329RrZI60Pr7
Wp/15mFq9XYmfnmkr9CKNoO5aG9UVS8JMdIc60pr06JfONjMsvQ8MujAmtIKcJDnd0uXztT/hDKp
69oHZCbIFKRfcbEAr1judn5kUK61/QNB3+twlNzaagbPfpPn1K4Ot69BkAnurveMWwNmnI3yEKQk
WKXKxTuHb+rBseLP4UVdVugLl7RsTV7SMiVRilwckMi8i6lr77ScqLxyNCKnMeaV8SukSVu0tt4P
S/u+rIUUZpNLkhvTMwmqE5rxN25M0tKyoK6T56MPH20Nn1/iViz8eYiXD9Pw1HxkvE72tS+r7jn6
ORe2+DZehcpYAxYZcWQR3J2/l8We4XM+u83BX1qvOiCe3oGwQXKkeoFLVRaXELxZmACtlYI3LAVv
2BYsxl77H4jj1Hlk5WkmOSCP7LihDAGHrw0yEYf9Vsw10hAM0AuJ+lQaWplSO+t/AewSxLuz/J2i
WsTQxxJfcqXyRNgviqxiNGyhtotH6KTja2QLzZFzIFxcj56/8KZYkmgiPOt2KcUqOjFpHcW43vYG
crdExSDLB488gI8k3bixYgVujpu54qCZr86ysGqUyoff+MXDCkiCMl0ERoAVukuZOg31et/+Gp0W
zNsmXBNHRysophrTkndgdTJz/k8QOMPrdQbPHJCaGJ73ePZacZF8kPJjig00b3qADUewocu/UUoL
GQ8rG+m5TFayks+EniF0LwPoKv0OXLsd/mg+6DGaB/GurlxZ4SGgYy/LfaCQKpM2MsptXCKRaQPY
z3CshbyNpLJ2ReIh3HLr26I1IDoqKOh6v6zlYeIwIJ9KTqvaZfkvcuMsREvkl6B+H14LObyiCyYa
GeM/d13WkQadIPYnQVWQVbXfC81vF0bG/T2+dJM4FtsogYQLtTeX7NRut2bm+BX5Y69+kAPFo/Pd
sVMQda+Y5XLQWG804zAI5R/FWxRrsBXVdHg5NsAyfBWG9f3wOL8AXF0oJzrFH1jdGvGBMAM8oBnP
hWr+pmq6wSkPf+nD+RXKXjhpOtVSB1TaJLe5exLFoxX4kC6yP0pPOjK2/LbprgpfPuHrNDI+7fLF
mgxcVH3zvbF1DmcW3djjbnykQ+rsBKKlXqjtX2Hr6xS8KyiIYGU5Kp04dQhw81qnNWqELcUT2sgE
awZra2GusP8VGIbNycfmF9LD9WWGjPPBlT1fI84k9Fws06WbqkkptiSmtEWnjhHMGV47j1DW3fdc
6KtG7gMchoXvyp7j3ESpocu3Wn81W5K+1E5lHw3qA4viQY27iOVNPiZpeKXVCuyDtLj3lc5nOBNx
XBLDdq6sumeT5PZ+cEfhnfKx4/8CSwlZG8FSPHhL5ku0rmg4D/6qTy5xx9I89UoflEkwpprTk/85
TKvx5sEVwu2wvtl4DVIwbCksl4LR+nZzHPQEOxHUh2cNjGlKMLrs8VcBjWCuwhG+0PqxmhotA6Iq
8qBURN/naplnwMiRvuz5nN56+NHeGA2oM7h+hl/p8FvsbeMpWzzPoTYvdHZ8m3DOQ35b6UM7KNZ/
ieEuQO7PkT/JpaWz5sNgLBNOfpTGqO3W47lqE1rXsL/Bwt0J4DnFvz/OOHrW0sxNWbnC0Wr1YlfI
mL/+5/VTqn8b7t6XcuitroN7z9x7pLfTukuwZGjlfVbffqITLHk7Fbn+35bn19KOnsy9FvhXKyDE
lsg4l9EJTEDywZ5RHhaz7fFkHzphpyCjwkAoI+SuF2wZiksl7gZKC64+Jsmih49366T6gUbeCsDw
Qxm1TWkxYWRF+mdaiJx7KyG2F+Pf5jTou4ChHaM5UlfacyYMmACzqjiDaNFsa2npiaIE8nPELint
PX4YoOaSOZgEtavtCSgM75KX1CcwRkeXrYsB3oqo+O86NrEnXwMahWJrLTa3ZvWLzL7cyWRaO/PC
CmQ3UGwTVw/PX3j8DV6vCjMTVqiPNqO5Ur+2i99Y8qVC8vLnFcHLvq4A/kTqThNiwbifgjb5EBZs
CiLZj15/6JnbNoM7pZM4TwB1kfClAMWihlEGHRJmtWIyD40Yb7w0TL4nDn/oYiqZnTFtytDyAjaS
yDNBCUXCXvSJNOBA8z1IJwXC+XGZrkmKCindTcMfSwlov92QvmKLZkDN9BsmtWLtZKRnBXX1u/ap
NWn5K/clVN2e2BSXEj3HHfnAP3PsHaWpvgZJnMX7mcPyMSBq7vTuUWKAMFBhu4vkdFZKvdiRAPYU
zjVU04n9WccrkMgJD6FdZdUp6aY987afkK8w1ARNZblq4cFYHsJN4EDM31nNActTIm4xjSYNdWoN
q4WooNr/WXAbaolIc2J5EdWMAPXGz6HwGoFvel5d8c+Nwz7Xm4AZqj6MK2XnXE0heb3xMSNXk+m1
BD8rJXiN4DYWaDop/4BqIVxL1GbBxN2uNLJ5vG7yOyZOqGAmem4mmmqwTTj54uYhU5WO5EBK1xG7
ZC4/wKk1kmQ4sqk7Srt220NAsk2y+tBCsQlY7DD4wzh4pOT+y7sDnYY+fKtBa33+1ccAznjKE3pD
ILCHJjFfLQc+tGp3Eju7bRH0pOsjhiPCZoN/apiXjDxByik1seuZ2IdH6iQaZdYdFPrwBbw4Zgjm
GQpkr8VhWER+HPW7MhQS8HTFU3Tx9paQfcoIez/hl/FekHU2jI7/MZ1RKvKDalWGAe1AXLdLTLck
WQIOEdLk8fl0Dfo7tQyi/eBkWJpMFIdvQubBKDHqPjltMJg+pwL/i9fFiI6GBfXyndpAKPEyA2xB
tr5WWXS74OMdf6MnBBdGqmZKW5mzS8CW9UeXQq0496XObzaZGauR+9PfgK/w/A4AWocAgSUVHNnL
rcvaWcTLQlUB1Q6bwPgQJx7FPUg/WxixTF72d2heTMDzaF/5deHCaDVCf/PF0ZD5rtmZzGmHYKEd
NhFNTsoLm91e7LLczz9zx44SqdCSciXVdqjIIxtx+ZM+1A5jIKQ7WA6DzbrZK4SHYA1Gy3xvlQMe
6zxWI7KabrjVECC+uTPMZvKkXMYCZk0JuRjvbE6iDyMzMtNONteec+IC9U6xXmF+X7LDEAg8wC2A
9DGnGHm8GRP3WXXdRzOCYwS7t1MiutTjwhIRSK0cIkJYKCxofKgCAnMGwHgcRpt1MHG2PE/YbTOm
RCD1wu85nlNEPc8l+1/2H/jHQFlnti8iHJUw2kbZ/f3xq5kdkeS5HarNjy+I1PqvyMgQLHBf4Vfu
K4uSWXzSuoCS6i2ybj+3PqRAZID3BoUcP+ikqjckxYNcmjaFpx7dMwRmOhhQQOpkPzQUu0g3mi/m
KZOkC83uXcpgXAuSo1pcUCLMsGV5CK2raSQ40e+oaahJBfPHNh5dhoL/CPJb58daC4qdKAi4n0L4
gQAq4EFaIE0HDRuQEI9LVmNeY6pGcin+w8c8VwqRkv6PsieHXBjKsZKzec4OvDTaIrXtlfjgHCCN
GGTWDMGw6VaBenUh58aTWfmD+aIrhRp9P3oL/s7Xlv/gvz9CRdcM++xCqFFEDQmJno3ApzvXvKPu
4w+/MazGtqlhc+3jr2580NA4E1GVT6toDZ3dRmyOKfj8KY8b6Q729zztUghMAC6SGD/I+wBXX1NH
lRWREDhtAX7iTVE8cyNkm4Dxmb4RK4wcNRp7USXjp07cznvFGWh/PHsFdwSgOxfQcsSfSWN0ejIH
7d+N0ahjUD7ZhbP/WRJ+gc7AiwAHi9EUW9h79Qrx/RGfhy2MmFdajeCLV2e/SgrDvQBi7022/ViO
AXle3F5v8Fkh2ye2bB9Fkf8ztS7h/pxAMJ4hEROjZWmQf5u6lpVdE52FbmM4BofFuc4dZhkw+zJJ
sthepMqy5R+ko/tyEwTnYLSABO4zzR62On4tf4ekHSz3MdpqQxPU+89/2utiRRjGIcOId/X3vKOx
8wTFmRy7NJ6cKeQHlqVfBor63V7mF8a9f0H+NP2eacm+1JuAoAdhfOervcOszC8AlCeQXLBUmZb2
tvnz8swygP/YGFhKoo/bVx+tLKMbNhHaCzbIx5HgNoKbIWgTkOypjUK/3y+G2SxAgwqeRdvxIJDr
T6SccXIXNj5XyLHu9+HnomnE2a8Tr93pLDQt879DSg5KwzZXnyLGLZAJcc2TKPM0XhmTIY541xhy
9Fy8KPCNk41Xovh3Q00UfcD86lsL0mhKUkB/GtJ0SyEsHG4cH2N+nuGv1qeNf1Uyxd4Qe1wmMSCa
F/P8PfJicufz3IC8Zi7q9oiksWWdiUT/Jts+aLcKfF5ZB2QqQudGoRgODGfV6eTlSP4mqHu5R53l
ok/grqwjdMMtjRCegjsrsNubluck5UC/sjAguuPR5nb8cNjzeMQkMbowchX6W0criWJXzpPQIglM
AIc2LvDieU8s5SZtXNvlOx6Ki1uwcANXtOMvn3/k6oY+awgVMspvQfGMuiz5veIaz1Pg89zro4T6
gAPepikLaiztKyrUYGzPK7OSZk62W7s1ulP4K22MH31lzryAm1CvKUL3hZ2ewGo7nFif3SuGWHWa
wG8uqVjhlERcJll54mS8AARHMz6BO4zBkNz77UR/iWCTmYx1O0WS600mTM03S4nZcmaUKse5/F1H
VzaVgqwu+BXz3oKF47CusZ1zY1ShFd5ExqFuzQNno/CQgMwoaI94bmYIlcVDrXK8yFOuk0sc4E+s
8oNcAXJJN6YACpaRB5dbPz23zWyF5kT97eLtSQonSiddeD++6JhRjypg4hVNfSk2CpYcm3aUlDkL
wbxyGMwNtiBuJAZjzjtiJRwxcKtZZkSUwaFOoBw/nrZXMsKU9Rc+rJXtwo37+qVpUgmNNZg/vKM1
IGJRbV5O3umuCnewr7Fu4WCyU6h0J1hKpEwnpCEirP0wm6zH25uOOrxuKMKVJZOCTZ99oBueBEuh
iZJaYQhWMCL/to7yvPA6Df08dd8dmOhRxwk1Yf2Tnd13cHrwnvr5YW2C1b7cxHFTCJnzkRd2mdg8
IpfsJNVaAOAXFjpbzdxDr0TJyaFVwVXUDnB6hGVtcMvSesIkutIHJ3oz+CDU4k8x+fj/97Q9Iyc+
AcqrBl1k4StWFq0BdEBokVFsRPQrxDel9vcoF4L5mYsEANgqYVwb+I1QthC4mtyBnAAjIa74W6xh
d4XwEn698DvfooQ6cyOKW9dzY1EWRkBXfT/Hz1MN2nzwSJ+yg2nTErIkzYsQaR8edzjBN8fd4Knr
2grb9aEhV2j57FmBDhyQfoU3RoaWlJsQsiAhr0EY1ju0og6en04ld3t1Tz6gbmotZkJxWggzIhVm
iTicXIErRIaxJK072ZYSO53IjiOr4x32QYR8dL94ygzCUn5CkBNO4J9tyTM7UaQpV2dCKUcPEcZI
pzVw1pPPI9a8bmYJGCmNw5AB8bY4RNNPvWQXxWE+AdxJCYvjcFYdjq1uaWo/sia4+29XUva2I1U9
BfL/Lfkrx4PTDs3jujWDLwFLzpztCoGK0F6Ue/PLsHkRLieGazp8Z6a/1UyES+xSkdFz1pz129fn
wFhRHACYJBxBQkqoCuoQGvn1fgwZXff46+fS6upremS/w4gQruiUBDZXPMMydUJnqMQtzG8lKZta
85tV81fAHGOTXw/NDabpkGTUfyYJI3+3WDzHKlmXhPimf5NdEGtdmx8ZXI2/0sLyu1tCNLnYtm6d
z9Es3+PHdIjH6kSPqDZmK9UcPWkTWjvHkCrnQbEp42MXjOx6xNQ9RpalhYW4MTjQBL4XY0F0rN6W
6figN9d6GmEHgxtaWw2JQ9uzy28Dp6KlRMEeBmYi140LpjSiKwAcUgwqkzIueRC2F0yvWDUK2Tt+
GHZo3+SBXFyI32N1qF/VJ8OkXj4ChDnfpJsZHQChGFKzKwKI6a+ozYsCRn31CXc2SEbb4e+RJOpl
7CZAkAb8dVljUX6fq+azJznbuvG2lfSmHuNZePwnvLl9Li11xhRufmAYK1dU69EmskZpQ3Q+2XZz
uqRxyX6qOmu9kg7rqvAv+5hwikqIGLtxRN43+NAP0Xvb0x0boEQ5d8CnbnoyrSsa+Od34dpUeBzq
uXb9cmOVARygxy0rmRHL+n0heLsx23QjTdReC+EjDyQW8XbeT2KFsGVMMqUS/FzczCx7TsFEM7gT
XzD0i/tKXe1L6ZNGrHQObDPtQvsMMxXCsFc0lKWY5lzHoYxOsA3nUFqxKG16ZPbd/XqB0YnvfKA7
hY+0JI5DsvUSkjQm0Imesa1S0HL6/+Kw9Im6wsAAU8A0pmERZm3sYFr5cdUtPBeHlAF9OhRQhQ/u
uO12KycOlrFYPbKGMuFea6j8UdsQI9AOZuU89Uj55LeM7JqXXBBYEYiTJDLV2jC4UpEtdf27hwhr
scW6a54YuLj0oUdYZyx8N5IOouvoB+yIkyWQFsh+7QTAcrJngkYkHWHfN2dYVB2t7fydvkTWst5e
jlswraZ+i3KLPAVW5uLCHWxGb1LYMeZEBaEsDppL8vq0hVuVILTGB0YuRroA0UM2AFtlisTEhtpj
R5Qhmwqp/9BqFIh7+lzTrh6EW37qjGOjwvFilrggTGDN+cTkQSNUuo61LCmMRvXhkgoO7Idy9gxC
a9g2qsTPYsrHXam7sDw5zcoIP5Q/ImTRlErph8VoOoAoWXAIK1ZkofCoYFu7q6oP52OzgSFBvZSz
n9VHco8NQGI3S654P3dBOXWWlbZbkXQ63M5j+0gJVyK/XNRA0xHJXJulcfi8dcMZ51fYar/n7Lf2
XFdgK31iPPiyT6CncuYlKRTT2XjZ31nA0+8c+liCTXYb/NixgaTXCOa2Y05COKh2FEtzzJio3vVN
xY2+wr1mxEd75wNNv+dwEGTugANJDh2bCwy4+jTWDdcsJJ2bsdYU6KooL1NaaChBWTh72Y3p6LxK
Y/6brTYQnyKRcNYZLl8cskxGb9JevPYxZuG2sMvWebvq0Ng1TK08T6vBsumVOYO9XnfyUn2wee5f
nKZPnG82X6SoF9E50hhWt72o/iCBCYX2ouz+Vc+Lo6GmPzuiamvAFMNIz6ZZhzJzbrTU3W7lZ0Db
Mvu28wQW+nG84X+Ke1AFLvN9MP9jnis2h6mJNFDjtjBmNbqFt3YQtSmP3+ob0L9ee+VlXI44uVst
GK/dmFJZFhsujdhs1Ab/HHY6yf+u2OA6G510JUwDQ1Y1RH/xS8aiOSCF+WEiCuN1IlbvOWm9BfUI
VsaSTDEG7aIQMsrPAq6vsUg4oknNS16qTdK8k2V4P8PAefO7Am7xly5wRM9mxUtIPeUIFS8tyhfO
miR5XSw3giwzNlia3rBjA9tGrASG56Cv5qQEZIzf+xI0s0KS8EcOb6yx84W+yD6Y0PQFSRuMLInf
kJxs6KUFm5mb44uRJzwgJMMKfXSMvYkFLHBjSGzNnwoxnliSCS660o/Lom15sWc23ySI7TCj9aRa
GY4Sr1H4OJ7TFsT4UaymF1RDD3v/kqL1JIN2iayigM38DntGMqNQJhKC969ZR2NS1E4+HhOYzIep
06Sdzh4DJdi/vexpwsHocnrXMHJj6+3ehEXD0MkNDBJEFbYU/pxCsDBk9k/4pxl6wMsOyG1G79Dq
Z+EFp0zL9v4BkKsD10GJTLQ2sQc5DWhWmbY0Hto16E84QSd8on0tHAtu2KQqp+LSPtO7RxqJJq1B
rFH4Ujk+vvSIhgaezmaBCDyIudvZ0A+a+ApkToxgre3UZ1RxdryiBAxkj2erXogFPsHbXzH95GFZ
nK6iBXAkVIMswQevIzmWMYIgsa1svm8m8mg/L24w272meN1Hg1rdrcqlJ00d4/jsVX61Zzxd2TqP
H8xWrP8Cn+q7xJCN3iPx84PC6QTuPQVMIod2l0dEyIqX6/dFQ7Z+sH8fJggT0ZHigvZuz+S21Wwx
LbHb1+/GFIS/pViEDEtlRpN32yB5fR5CgeLHhq2lcS6VgC7gbqgjjIvxYNT+TcoWWINkyadbhmd2
CIRUweD+OEPcouSpLGKPH1KLJvGKgotJVXXbYsEgzMwkoCKCnsxh7GqSsxOq/iq6rsd/PjK95oIy
g2+8UeelYS4xrMWlchDFiIsGhcCbeJgus4yg9e3PidD4nypHJa+nZ868h8qfbK8te59Ml7o5fmZR
93bOH2lxaXFZREGE+3twT1fnrN75P+7kF7Xr0RmX26S0p8kEaMJeFfmW63yexgoDLkdPf0HFGCrg
KBRED2SIGLSsVAoNmcLOxTg82hycZ+Xf0A/laix8+NGSBxIOarSFF6rp0GudZKkxG9N17QieT/U2
2rPFwIcpwC45d9Yt0RL3OkC8mE0AgdehPYjsHrYC+kK4GN4+c2SnItMAtLrPhozXkI1Uzn8TNxaJ
9KIKLWtLa8lf8BUou4zal8SqMFH1frkf8uyZnEfIf6MaO4PM3phPKcdJQzvJ2ZuxzQC9DIR06XGY
cgsxcmnv+lPIH1jvD3+F/G2lB/UjKHbniH0LwdBqQ5AcYSexmbhXHCpOPLGsJh3gVXVeHWUNZ8XA
mQbvROgTg0jeBKmEpNVEyxtcMqz21NXjZXxjzI2p1ss48MPDg4a0WLlzYxVknP9lyMSJ9CI0hNli
qSsiCwxV6W2zm2yBiYuZrQoxLr6lAAtE2m0Yynt4muZHU3ORK4yIbeASUI3eAGhESrWiWS70oGPR
MipPfVk16pW3aSiXFVFgOxF8GqYJ1gD4YeWdQ63SPpvIy80fXbIAr+2OeXWIZL1cNLkax7vvKFsN
zlGX/ZR5XnoMjD+FCTaUENxmDgJ/M15pbDX5JKuRBY3wJKGN9ESZAX84p57umd/siZDhy+PYSiIi
IZa5HPcr9HX6jjem8LvvFLTUnlSEkLVJgygLqR54klDL7ljIadidW2/KmkuD+p1KicxnuR1D9jXW
19uMNoopkSQTFAB7diSIF1rlo+FNXRPI/3u1jMmlfrXT03wbK/CvY8qIVm+32p7uqKOYfchG3Ko4
hCsjT559r6XsYOmlUjMvwrqB3R/L8snABegso4tpBx1RZRtMtgaKuajp61PvKX02O/tbcNe6izXv
ZJCHFuJuKc5hxBXTiENuotJbEK6geZnYB99JKpBgG6Mo25rILmtJXfG8I4zVAEB6cmDa93XcegdB
aQQZrWGrVVpBLbHO7FacItOypuIKd9thxKSQrRSIzX9sL1hdPoxeHFSIikdsDs2BIQkyF4qzDmY2
W5ryO8AVB4ENLEECdnzzjzs05UJ0W25Qk4OT2cEvxlH/oT7a1EE80eaqT+Kp8o/7OFYuU8ObjA4H
XcTvHhlOEHPI/Lbm+UpCvF9ALRQXha3k+/bajmbX3EoLB/27j2WuV8LYYSvxN2jrekt5Ciwud3xq
eGP/rVuqX2ubnHOf97vuKrwQqM6E9JXO29bAVYMhiMfTKDaNcEry+14hkrku7piYudzlZaNAZMc4
2/oaJwqsxCHj7haTGGklEmvnOTVlx256WBP31DU7EJzS6Yn9p3ht7hTiOi7aFQidy/hMCSh15nCR
+9SEXrHAbuUcZ1qArgmneWBw2MEzqqnViZip2IKiPiMsSd4GuHxuyEfgCHxvWZJpGw7F87kkCG/E
muCNW9lW8zbK+/Z9HHIDfydKJH17ZM1G9xknnxsXaKz6hmpz3Ep1bQRON9qvxCVPDuBeAV68tcYS
kCan7GawKM5+KiX/tbiDet8vRsRjjtHs67hg2FtZHB6m0d1DSQzxYWVLjU+R6RXAs9RXGsWckldP
xGAxufTeh+iz2VG/zswciTXWjJEwrAl+kiiWL+elyBzHlGL/bKcCjSDcaPg7wx2OvpYv0B187afv
b1D2PDmrVTJm9c88PjcQ4y0P/rFIjVCb3WzxxHRu8BkC1Ts1osVyvbQ/MDxJ5AQm0dtHtAojx/rV
+rbBNYlGZYGgFvUEDAHsay6ne+MluV5w8JTrnFsBHki3JcHE+sqT07So0gH4HDS+2EUC+b5UOlKr
oZ8YMWWWDkNh/uUuNRVOIsLSBKNj6MN5hOB0NxWih1YDEOEo/pVwD1oEuXo1Zsip2H/CuqntlC14
3pSciHfDIzYMe6xmxPELXj0HPqOtDfJgSQBqBWkq9VndZmmYhZ8PPLW6AWM+RbRp1SL2om6tR0ZL
QT1fvGB8+b7cPFU9VukuuBmsbupQU0225f6ED89Uv011sDQdITe9boajLyH1uQvwfIagLflcmorO
yVLSc6OTsUq0NDrG8h3kgI+UWCz+usqUTQK+poBQ3CSxISSUpmrrhI0qdthvAdzqJzUwyUiYyYb9
HY+9lpDv1Jeb0dyNlGVvVIYsf3B75xJ4LZtDCZegH5G+dHjl2knh3+3LmlqNVaHFerTvH6TGDpqz
bl3XQpEn8bN11F74FHuZkWP971qeQFzyWzx6mkNVF5qNnOyQHa5AS6vLx61A0IQqkWWoQby+BJQU
lJgUfqKbTT65pXGnUJl/KD0GtnmweU0XJ+Q6yf8K3ibZvcj20o2NtTL+KkpIQE9OGsXg1+NN3wDR
sNR/SEoqzLDYa0lWP7OKWic21JWdw1Dv7RAJLXH6i5XlSxtrKQtXn9zJHECe2QCd8WvqetHBkzMD
Ei+AVAkOvWRZhRT7fp+gKEwm6o1gF3KfKyujtQrdfAxZMyUuzS473l3wDHt/NairKCkOEj4e9zhS
57gHtg66CGD5vG0SlCbpv0pxNdXPLKo/dkwNPvd7G5oS66jcvLT4cYpXV2kZ4t7RvzAPEY/y2tr5
8kvwQtjQosFxVus53SAGEFI/NHatR+wXyUOTWd1lxjXKmy03Jq/Zr5qbruAWByWnOiOxdp/UGGjD
bZkbZz5+H4u9VMShD+ShL6Ar2j4hneHqc/FkJYHdfCNTAjPtkruAyAHxNwDeDdoTXMhDMHULlWjW
q869Nna5BoU6OpvLWhKSLKYby00fRIsLgSqRjvpQ2siJFg3MYpZZDdoXNhhaku6F8NoOtIMRk1LC
8k4impDZSE2vsBIAB/qn9bIZcdJMBQZ53M1cgKfe+tnSw+1wbvE3AB3UnfnsWqDCZuQ6CH5NU8BN
6poL3GYY29eZVOocfPYyyWWgKDkNODeqZhbh6tqukxu8GmhFHgdHglcYox9J5YTUFxky/hS5RX5o
1KQXJ2Z1j3ZYNVDOU+KA/RnENcmCQ3wYKxjZr89CYMp47/HOoSfihmDKyMTYmQESBQ1g/Uf2CHEo
dUc28Yfv7Kg23NBVURfa3dgrVP3emh1Uq5F2pUtbetYbzCM2CWyIqiMD1yTuVgNoKacZPAKhtVWH
HLS3hhJG2UzO6qJeFBx7XZN8hIet1JAASTPG9OS7gC0PVw0pKD2KIr6KpqZc2OCJy2yN941817ZK
YGfF6S5FuXv4vXSoNz7P71LdAUd9H3cwfS2Npm/ot728V949RYWvmOeKFMXe5Pbyi7qfAC63qPNM
ZEBOWzwkH9VUAC9179TIQxI4XvDcUHlhBle2NraMW3cc40sV3dp4WwtLyTsmnltO/pEYO2bWdvuU
FI7E/7VFYAfyaTIouRCOEis7ZS/9sutR77qFz4vIyVlj6pNNwglnGgPjBKoqpuEhdUioZDW6g+zT
qdpDXnIK7xJ2546gJch5EbKfAF72Fjy8hPrQyRPrUZrHzCMm+io9lGS4IgXXzsbCzX2ZHD68OBPZ
a1rN5slb4HSuhzG1otPr/uv3zEmmZXX7z2KkxTzAV0wHgj082j8ZMrPZwMorP9SI1bzOQvy+VCPP
Rqn/dc+rLpzU2efS5HuklYmAlAVMFkaCed+p1hFg4/TH+pTv6ZiqlAjLKmoHvIo8o3WUxqSMpSuw
//L9o+kKy9I+bnGtDS49VfsEJNDeNmGRKyb+YMY/jA+eh5gLM8oHQ1yrBl+1iS1q7yHwVTa3hnpf
t+qPC7vQiBS9NiP/oLY7EszVWFUqTDr1MUE8cY7Bjnv7BZ35L5JJUD3gFauslD47ex4FWN/vHp88
UQfE1WaZ5stpUIYa0swo2Gxg/nykvI9Y2XMsQoF1VJmDLxlsF0dyWxKzirH8v85zdX49iPMvi/H0
6QYTFSTeMDiQcl8CCYebTNVk5OzXv/AsQfj5A6zPWwU3sU9CYNWZQKr8R8HHSUZmtRAz6NzhQPj1
08JyuHGHPcpjDrJivKuwqH2MvcGDSiA7l70/d2zuAC0hxj27ggOWuNJ5mLjYHJkioTsGVm/C4jAd
+tJ6d20T/Zz00jpTc2And6VqklgslSpsq7cahnA5ddHoqhgXCNjhF49FNgkzqxW6furJ93c+yoJB
dYVI66yNclomcAGIpnB+lzk0k0AUMa1vlNtdddMSl5cNel/rwbLK/FXEUcV5VWk+rqTBisTeEGMf
UlnWoi67S+V9OuAikrqHlbRTv1XLyufF0zO78jMgyXmgUNABEsX+Q4ujVQbZ0rLUR7JEPW6ijWcJ
+tyPKvIK910z0cCXd6I/qQAyglvAOB1VB77L2qlH0N5/5/K4qMVsqU7Iv697sw9PShRzcsNlxS0G
Vxnbe7kJremqefTqbYUjJkGpHxoMyTbSDIRJIMRT+SIx05euLdI1OCrfkTAWCu6n8S96mvESfV5N
nXGhzB/YRnczKPt5iKYuWQ1P98/XNBK+qvA4x44VgzrNgMM11hhTQMt5GX6+EGr8DQ1xIexmZsy9
WnZkGRBkqMF6VqEJfUZNR9wltyD4KqMSRz350BUVQMYC06IFDzBACNPaccxTLGjQK0ZmVi7pMgcX
b6E8DeFp0LZmhSSFazFK7QeOzpmM+sBQVvkjETRD74dkZR5krVnL6rC20aemqtiAIgRWN/rj4Nop
DtoJzfqqIu9BAuBmZ5u/wCQYAv8Dagb5OyqmmyisQfYtPHId58buXd9IWmvmRNbtHVOrx9Q5NhPB
d+ZNNf4p69tmwoGOdDE1fmHG4YzkVrmsnHoCrVtciDNfwx7z9VhOIiJv49uQNIHD4vll4TZVAPhn
SSLa/wJnxiWitmTERnZ9W6rqkOfTIDbyXDcT2ObTjQjeptW1HSz3+vrfB3MiaMRRFZ1g2cc6QxFm
s89XoB/TY/mJT1w40S+sr43labBVeRFAsT/deWxYfnRDzWU6oRP1WuuchVVvkjgVLPSRAaO0xXnh
gMtl6upuLXl9IA05DQ9E/6q5dvtZH/JyL+R9YEgF+V1kz0lplv6jFn1DGI4WrBIxW2B3eFQIYxnd
5y1Dn4CNCkRbrOgC4Z24ySpRVOszR7YvJMml/e2oCW4fcBErgOxUGsWB/eui34S4zHouj61ib4jN
pCBcYQ2acSItvHcBXszHpx8GsPYpMJExx/+73XxkR9W8wD3TXJq7ugoJvzJ8ngQ4zhwAV3RSKxQr
Z29gV9/QZdK4nAEawJf5TrWaY1id9WGU3pahED5SOw8CCscYsUymsocjSBkiGFvIx5GpbfeSDeSd
ocXrkuCxKQ2dgGuPml73WCJ/esAF6BL1TRXIdLHsc62lV7bQRQ0Bu3Lt7TWj+/t5UI9dwCTiuaS0
arXcojX6DfjiuRRgruCyq/hVwGhoYnoUGKqXfmkpH94bINEt9LyfqaEAKdzFff29qtrfWPldd3mo
LzXuSlL3d3Yr03Fbveg5sggBs4t06kt8UZWeIwVNOvnrEDe16RKGyhRtKt7zNgTjvGdPWIXCC0n/
oH5+aeuUg8aym0fwQNKypbISj1T8weQLqjbxejdNLAOpGNk7lfgE7PMQw2VFUdbdL2lQX8HypME2
XWJr9TVJzt3GWgNSEbdA88ioFwPmEhDLN+poqVxJ/8s2m9ZFQk2R86rbovwhVNWrNcAWHukvrCeh
yMnNqBbIgIvN2GU1kgZJPpKKURO1o6dkqQSECU9Doj6Wgn18oHO1UpIJ2EAfyWbMeewDCyKTn0oq
3Ew8JAJgmLGYRPQO3iAUpliV80CugViQ8qMb48ioc9Hzz7RhpN8l0kMeP/UByfu6P5SPF39Zlrdw
rHoxqZMle3JXtMHluuT8IQln1nIFQ8Hmbyp2902CcAWsOXq2dZm4M5Y5p4cVE0dT32i84VwAP5Gx
7J+vzeSTxl/dOoIMpQmD9t28FRWYKfqN6H/nOCC+fKx7SvV+7IFULuLh7pqBIEa6tLJVFTcb5f/F
GhA5OL2VO2M+gYR4yK2JokOkC5h7wmDGMgwGZsQzBqfPmYDxu/7jb7H6L0EjnBVtcbFWziq721B9
DMHp3QKETwFvyVgX1EcCGjmumcxFnggiGvFy39ZscinvOcYc0L8agcynT58bpQpLzJvJnobuypxS
iUdan0kO2kK3lZITGuSeYcYYrh2j31SvzIR5KL51HJH77DFOL7OP1l595qCrlAU6c5RG/VUz+LT+
jB5xHW11Tt6tzxdLoIJIa0TaTGOP7Z4ypEyxa6wWprA2sUWaz1eXBUfodMb6yqvGkUyO3r2NiPDQ
73qfKEck/hiuI66DY7/CThCApePg4fnvcGhALg8t/oR9tRI8EEi1D9REhOhr6Nu56Imm4MDqTCHb
JLJkGIVUspX8JgOS12eSD8yFLx+HPdI132OeBbkMI9m2QbYwS4wyW2IJO9uLvFtXh89oecCtLu9N
aIosb/qLwTRshP6N7ddDQXF1Z4oogxpz1Gw8JPjlYIMT9jIcm/mkU+d1SbQrt97s9YmfhHuzfEnp
CwwuD63Gvf2K/xqvW2OpPy6EmlNxkvyIfLZr75lbjsJfBE50GMaiwpqSu7mI/tEFmp3af9HRLbBB
hlL3v6FRyAmvih1EnXB6tVGxfpyZg9kgLH+I/M45FQZ9L7Nd6GlYciDRjzcOgNPQuRn6TKqCTuMx
SqTvosKmoXYv5Er+BYm8vs2seRNeQ6SQYI3dpUyoxmZj61uTl/nabyuLLlJWUHerkEpUEKq0SCbt
hvjlhY0BK4rKQfLMRa4BQvLV71RHqQckMlOrDEywIqd2BTUbg0fzO9uanKglU8UZYoEYyDzQUzz7
S1D6s7aMdex+ecF5L49unX3BsxVygdj32HmiVZ/qPBSYKCf8zQC9Au+3UA/qqPJ2A4vc3rUKT9Ja
TVIhGQkho4TdnpZJPtISImRj8xAWsXMlybUBZpuzaYRiHIRuJYrR+oxKh6t3gPp1C7xfFtnmZHlp
q/TH2iAtmldbanJkyx+aotr+oq7q6vJeoUCidvpvzh/JKAJaDtZpA+OILyyJ9of4+G4h00swKc97
4lIbRXGs31taSWI07KbRxPJnDjbuvltBN6FqzH+Ar1LgaXwPJe1sdfh62OOl8eFcoVjIjZH9xatM
+TJTU7j8DD0/jswdSBaXn+lFm2rRaejkUB3vLbSMfkQn8ANSmFJMv3GV9DlnY7vNPzYq3v1Ylcd5
ESX5FXobZqK/mB+IPRIx0Iwzxz5ZnCgaqKEVPsQR2J7AVuiLLtmXoRpo+xHG1dSAhEeG1rsO8mHI
gJn8a+oCv+QYa0eFHoAyY7zlP1j+m5I7yvOl2kn+2IGcoiS3O+my+4m3N1pMJRD31mUPBgg/UNKP
MplgPM6gTna+cTkPmjnKG5nEMjYbdYsaHrY7V2hq/o6qJ/g9Km6VSoFJ72DTaV8ZlfvHQoWb3wpq
x3mrfuhyGTl1YkQZk0VHaSuD8bnbHBbFsplhWzytZX6AfzxkZZZKdZo1gnSt79x/j5rgONeQy5zV
XmGvIZOuAeQ8lNUj5EsgqPaf+aihCdOlpq3Cqe/KwFbnfDWBRxg7Sf5sn844zb3tvOOSImXSrSbT
DgmVTfEqkyIweLJnCIltoPD/5j3XsdKk/oFqFZkT3y8F8BO2Ftb+0L3LioZrDRLOXaNAG9SGPknO
4Fh7rQH0ZSk1mkU9ScS4+H3TQZPS3xge5gemj1PEFTtNhTCpgAmVsmzSMgPEnqsSGn8fo1bdFjB8
mAXCC6k7pTsMuTAu7MzpblKjZl0s5toAGSpBezXXHyXv+CWGQfHMjaTh2xZf9l22zMq+jWk/5BgL
wIV6C0iQBQPr9H0GEeUtgD62N8DHynBmiVNLV7PwWkzPu44k2RorM2zXkhWEnrEVu/oEOdyN8YTX
KVBFRIuvXzG+nGXN10QREjBixgJ08riy1HLzQu78Ko5L59ciyUQ0esCxfndpgqq4zFj86BtTlsrb
aZp79R+X1shWl94Y6zUD/NmjUjAbYehf3WrL/cD6lCMsLQvPtafz5arutBe6iTfWtNK/4coH0k5g
Q03N+S4KeOTtMPfDpBeNMzL/5DAosh4nYnaE4K/1SN+a/qMKXLMflP6rGWAmE5L7S1a/uSLqJkKJ
J1xO70YCYfIaqiMLYDF51J98Wb4FRMzzmnPmuFXcdIjiN1veVbqX3AxcJaL/kDgs0f75uYGMM8e5
cXpR46K6CW+sjS4dio5orGy7HHympyI2Be0O4+CyNIouc6xJVKzfHrHZgfTMIx4uMU3/rBZuuTaq
XCO347PVtMaOr2f7rD2t8oQ07yBvM9/V2KCMy/TvHJMaefHCHnH7UuBErDoYg6yx5kK+vuQ5//zu
VQisEayrkGGclSkxb5Xvc8IBPTRlaknyx/hglisL/5U6NV0FzTR48d+j1DkSn6LpygznCHc5mHKs
h1nE7EiCI16QuXAzw4VSUdd8Wh6Ke6FGlngzVv4aizeLLnwJ/oWN0+zJ5+ILrbOr3MWPo9RWPhtB
rWRrWFo82erb2NmpCfZWCPEjwwH6Z/lCIgGTgBzAmAmViPfHrYijawzerOPyrnBqYm8hZpCmdMU8
K1uyXbDPWc9IraXO2LppiG13f/OotJZcf8Cij76eUySr1YSvczy0Gyk1BsP7rIfmirf2ZVhm0vrc
PJLxQcINK+u1UTBoJ81Fi3tpMjQ5MQKvPPBCfg3Gljv8C15Ge8GPZwKnl7VLj+A0xCW0kgnk2KFX
7217nbb1jMLFzvWUC7rK8LaNga+qUeDwsaCc/4r/MoFl19zhIuajtOObn3gTQyNjwc7soyHjIU2/
sFYLpOmOGFKufhx2FBUDvIbnVfY8ejwxMZMdyndb3A2G6K5ztbAmhEFDaN/jgrLsxoUJ9/f93Fq7
CllGCQU3JetYy+/dpE+bGaIJTPQoaKzFn/0T40IPMFLba8ZbJWX8DDHRZ3LbSZ/OgFZ2G704iIKd
g2l5Po/vmE4M58KOJoJrc3k/faEm75nd1yuihIVqDmWzb4Kri4WW0SsjTxqF8qqTBKJArdLVxcrz
U3j2hwUDxfzkhPRhf+tpu1adZwx3xWKLF2dWgW00XlzHQUEJFD00iJ+fuvPOzwVHHyXc2bOJ28rg
1Q+MBRNHpfDxuReLodKrxhE5eKI1UR63X/blOW1e65D0kSNSBiKC/GDiKRXaTk8ncyG6CtSv9RuF
QCBni/d4BTHGJnOLj7bLUJBhEN2RIZByLKRUU1yI4KaDoHNyHXCWCU3q/WSCP9VM+G28WcujCQjT
wYRadmereFGlMXqZmP2Jc86GxJZ8etyeD9iLJGdy4JkeuABNJTxNnzKPQKQpATnZIeRmjUZS6ThA
DkSXYsUk52XtemUWknHOVk0CIa3RUm7mMRxyx88ALhBjgIGvvEGNTHBy3W6KEn12Ug93yVHl4G9T
CZ7OSSP6mVoqc79CeZ32ioDgFDglUrEHfEoNc6wnMrOdAKD03tN3OOl4Khbfeqniak96NmlqnldU
SMOO8gCgZw1a3btoWKuaEAZx0Bl7vU7UfBfiZcd7EbVOSP7evv9uMLAGz04icyr7uzEj7eO6t3/4
R5KaP+m1HSV81XZB4jj21ZiNR4NHGtnABbTPTL5je67y91J+lhOoWsqiv5fpcWqsaMd2ag4aivnb
C53YmEqI7GnVirTFfj8PTq+7/Q7ibx9GUOd+mAs8ky3Q5FsjrpiYQHS6ixSGTSts6nsx0rhJ014a
TpJqpDracuNCv6A8ToiuYtlNy/Xx/FS5d7WUak1BFTZZPU1vGPHtp0HKGAJrBTvFihy9Zl/3/Nis
QRjkwswBZa49/KL0/TG2oA+LiMdBrOA9Lr3H2TgqjNfhFn/IRdZZXVQyRd3o/btfq65cvTiGfSuy
qmkHstGACoqsVDo+zIH2b8ly03v75ivVFvZTHuRkPsmKDPu4PdGAEwWV0D+M5DtDaLqLV/SLCrmV
ba7Z0yvK7dbGP3fjCTQON4uhoQU+ImHCHp5z1F1+05tR3jyyGyegiMql/ej854Yzmpkkg57EVmdj
iRIyZl5vMzcObe+4MivJeAQkC1ONilrfWchg3cxoyY5UkP8fAZMlWaofaHJJBGXmcsm0ggPSS2Fi
MeDaOr1LmdoItLni8dNgSWo6ouyonixmpArjeVkhuu19py7W6HLYQmko4um6tDkGgOJ52EMvA4zw
ziqym/RFIHRDvnXoBc46VQHdfYISoDqAjmkiZdtjQw+ffK4bbBQHoTu3h3oaTmAPFPEtMJ+xg2Mz
tWz00mO5P0v3HDmSIt3Z41SD4yT3vaMEkNoqRyn7Cz2ZIQwJUUeSGL9ImJXzPLZ0byfJfA6Zz3Rk
j96kNZ9iCVlr1fmPcwcLuzkXpfOEOoslST0YTY8ax18onfecamIZpevhPm4euNBFUj2uuEIBBbiH
DKaYgA66P37r0r6CdrzyXw1IpXIBhKuKGhDMcesPK92hkpVzCy0mceBjtVMtpyGdfg44zBBJqJGz
kv0YF2N9Hp382x44wr/U1jf0sKf1bxw8a/mKxKrug18LPPKUHjJtRoVF9FaBYVr9FRQKew7yFcgf
LyDSvf+EdyK1p54tVLOdwx8EFu5n5T4PNc/XJzjyOklb0PPHYdmycUW6TxWbszjDu/XqIKXzEup6
A0fLLD+P4e1/gNfvmzyVcjcU7IUVzXmZZa8oMgtKjWL1wVO9CIx4hK8y8j9HfN4IXlrxVle2N0au
AdB6zLp0TPfKwJamsXleVV9qLxnZztEiyQHraknQAwOXysyuCnt62MpXzaKVKIThm2ZG4v6WVmMt
UkHSnTdEWsRZGyrIrVtWSQY5CZjxYG+e2Cq40fFs6XIK1uW5vBJn9sP479dD8Ovv2NVQ4FKZ5+cV
HG1Q+OrhbQypxsE/IvyR0tk0bsGOODlyaYhpOJNwv3oN9PGjENX2eFOYN+pOFWDBT9JF29IwfbAF
msWBdxfI+IzkwdmE67rOCy9LAeSGmI/UVLPenbWvCMhdrqwKgq6a11du1C/kCugFwg6cc4HmSMFA
3eZ9SanXP59G1WewsuX/AIa2iplD3lU6+zsb+0jfsYzxN09lFUzgAzCl1SdiXQ3X2DTqvxq4EtGp
s136bI10jnlnA3RzIoSdxeSeq8BiOL6o4lp/1q45TnqZmCMrAhHZo2KTMMkeQ5VJFhydaYJ+fNT2
n2qzvgooXQ+tejAKA6SIkBGNzCFxmipVhQHCHKwlLk3fdmwS8730rZyOZ2sWYpQEvGG/DUxANTDa
i4eWTwQp2s5A1D7hEAl9T42pHSm3yCJCxoye47VYpdJYxCocgqcEzpozkbK3uUrhpu7b4MklirFj
uZhq2DUVCnT/1PHOf2L9HQO550es9A3KZTfA6n9jbkW0EugE+CnViNlnkyro9R5LXmMEmeNxFHtZ
Obv2VO5JqZQMwwYErjZdvYH/asP/sCzq/vDv1zitPnZzRj//7dDALmKnJnRUGSg6iyw3TU5Zi6YV
et+rjja1FbLdLh/EKnMAIjmOO2vAueUVRVyt9PMp3V/23I07h9rfp1zm0RpBmHuUkfDYUefioAc0
zxPUDt/LCduc9gdL7xMhwX+UAjpoLPmBCBvQiezXpZzZnbui7BdGDSQ9fUEOGh/UfKHWlz9zf/kF
alkv9+QOYtaRxHNCc9dOPn+MVIjUEzy9wVGakXT56zWqqnXzuail/8/2KHm37+S+e1rCmR1hkkFn
LtWcXTDxve8nDf1uIHwppWej44UjtDlF7HttDc6wRLPLkvHSa4nuTYjTOF0r6IKe51+/RZhd7mLz
voQTJfQUv84TqzFbaNmAxIskYs6MrqYJPqqUtZUDPvvQAhZPSESg1n+MAz8tMiQdlZgGy2auY8yX
XFNQYS7pQfv2LQOmscb6q4rWeYDVlet48qStGn7I3w2RjSejgqC/+wy59KUcpSzUiC8wxUCtq7l2
wVg6BDKiLfkEWkOp8kBOPpFKIvXJC/y/O2yUPwLX5m1IBvvo3SoppCcl1uZUWJBh49uXFNOpr9Tn
Ta+sOxqupbMEqmtgA0K4TbRB/d42FBGubEzBLbjZIbdJevUYOiS6ZCuhpr7amgEBrQ7p/5+uFRez
y7JYw4gyDbfDc90YRPrqgb2Xiwkx1ymOykT+F7C2HvuwHv2IDGJyW0+DIfYEZv+IgsYLSfNs5yFH
42CT62mTGlD1zBRmRZT/aOXuwBtyP8CP0PfwrR6Qe0fK9xNi/9UrMU2iRaJNPZ8t0yr3qdK28SQm
6VufBCzS4tvCjHydwyEUlHQZeyvvxnZNykp9KbM2hIELTXKYlbKNZ+mNL6FKSRO44o2H5jEc7n5H
5/NH4myZrorPs8dyd3wrBFljB8YGEluQo4Gb/Tsq3rVYqDB2BAN6D4JKLMA9z2HiJhgqZ39efUzL
nUcxjDkzviBU9gQ/VDGS7/rn4kR981ui5Mcz+a795h1idOQrm6btr+HkrSrb3ShkegGYh5bsYDTx
g2Lh/3bVCcByRTUqDaStFH5U6FKVCtVIFfl2c5gwPuMmmSL2vi4GAXhfWvuJoao/esq4GdPFQoDf
9lDvmfjc1/UfBzXnrkdN3HJ/h54vl+YvmrWog1iNsLm0rF3PR0AL7a38R9hdHWrXS2azwd+Ov3X9
DJQplNWhlJt5qv24mjmKdC3LyKkpVA4xTzeMq1zFM2A6PNph8KFcmMLNm44x/IHBqeSV+FOq/KOr
aNj+egOJhO2smAL8XmQtYQauxlWjRD2d8EkRs9+6NZ3DCxS8i8T/BGSkoR+kQbxgzrKBZXre5HWX
lK54JWIpsR7Y4OKwnibz3dL2ieSmnmhXTwBwVM3Axrn4/jkTuplylHDZlH+WXRhA3ZzSoUFbOELE
nvzcDUyRe/JoJWZ0gIPiQ63DAfHuPLUUkBi6xu6J0n767Er7v875HiHpWmmDDGYOFYP4fpiBoVSC
CHOKv9+gq0s8MJsLGFnqiJsTAkSyeQHZjsyIapkIdaOCjKvmxBGIvASbHyJ8GMVLZ6QEuXEpAP/q
9KKsF1cykVeUZtCPiZ/m9NotbEXF1jPg43Z5ifX2vLlpN3vNwY3kYPk/xMf142SJc4N4rUh/fVUR
bU+zpenz6mNLzne6mdvkiqaSKzb0/KrJfSwjQBhsdlFc2lcOrgrGkx0PWjX1wk+DRLsdvsE2Ax90
In4TwdgTBAzixlgjIkIGJ4S5knIXpTMHD1HCvlstuppPO1ix8WAXdnu2zImJn8XOFjugT/6HeE3C
hMVJTuk4zKLjJx3lRQRyWLGKea34U0SCs/z4KLp3BhG+9NGPuFDdKnPoZkfq3zsoBFrrBq+LqDCd
4ofrZMaUDra/Me00+pkF1eZttDne51Jw3alDndUjUJwzSVq4V58cVYeYKsvSg+38VXx+FaNDiROd
Je3xMqvtq7ewasD601eFFyll9r69HXKs2KO+lVg9GP3qrdBTMb9kxKSY0ZiAHjA9C/kqBkwCZ6B+
8xVbt1NIP6dl0Q9cjB2DQBU2UfPJ9XjFTVsEfU26hIVrTgsRVvt338sCRLcjZb+jgfkd0A4V1N7V
tc9OPQ89P61oGteaeTILSx22O5sqzUws0PazsUJ2SsESJ+vJg8NU/W4zvCSK/rO5kpaGfpsQr4z3
h6Fgea3KZk9ko4JgrK06rOehypCCPGO48UFxwfXJ32jU6eEq4XN2aJRd9v1BsDeneOhbaw+Dn3mD
1AsjjvG/cICXYkRsS4FMfXiY9a//7Rca7faLcvvCw5fJkKwyn6HvhPSQqPtIC8LlQFzghij63I/l
2RaIukzYfGjRO6BKGoY1J4oeZKdlh1AqJs+8H9wN3J/Uf0YJmc4NVkRQL6QPGn8EVFJ40ICxnbo8
DCN0ktQ40dQpYblw7r8w4YVdn7SN66AGIptZEu8AgbMnsQTDC2pr3HE/gCFkbIbU6hsJy1gs4rwH
tI1cBBC0ZUxZj0njwFVpcka1IFNX/VjC7VKOBX6LuQ6EncDS4rOzLtIwePYZ8RF59lR0VqK9jD12
vKJ8bfmLY4X7U/STbUbfErDphhJ9BGYLG6RVdZJcKann+LTGPAhtl0qVXczt21qhwVOnOQCU1Pvj
CgObVM+Tm6yRg2inv0tMA2RJoCXGAaX5bXCqv3WWznTF5N/hFTZou6bO/8tqL7zy0eaC/+UGBq5j
iMluJfUi7ZtbT9Xo4VoMfBlwO1U6AwqMI27rlxin8aoE4wZ4ptxyKCXpsbzqcA10r/sdBBy5te8H
IL5Njh77abHy11vKHASmZ6JGsRzcxu0FdyqLGmMwBbVlQJuWqP0fchWuF+5ziKnpDyJNEENxbqYW
2dGhTm92/BCcEApFzFfF3yBPWwFGy9f5zSvDG6P1vjM2cbYTw2GdYx7QMQtEubrmzOpcU9izo65T
1WvW3CML8GKXletLUWJCW0wodqdSkU31pst90mlQOY6kJKu4zu6AbpRmA4bqlEgjz+dlblpBThKY
oJojuijvi9+s7X4Bb6tZAGNAmUjZ9EtR9/Pn86HzQlABvSi7UvEZ3zUhYQD9I68orQfwAZkVVNRX
cN3R8zp9nGiK95JH3UXVcA1BCv9FHvHRq2fqZPMfNCnMCT2bPE+7pEEnVJ01Hiw+LCDesT7db92w
1XXBFISJFjyAs8KQF7NUH5ttVXC4qtT+j1el/FspKqV9wzAfRIPwNZMfX7z6w9BETmVRZSzlK/Zp
CetHFkg8vG/6J0Ic818TGlb06qvRfm8d+qXHD8hs8PBtfGjgyu+A/cA9o6VI5XKWomb3pTGhAab+
FiJgEHTpiLI6XQ33SWVbGYZxctIcy28ABheYmGq7kEtX4Sa5/NuyM2uxZBU5hszDBGso8GY7pk8r
tDPxdZEsklmOyFO2tXkPQ9007KZGv3jckJhtC8HM5LsO/v+Y3vGJ8NL8cmI2XQHASBVOPtVV9GFN
FS1WNZUs9raMe6RVCCO/oJqnD7qJtyD8nToy6tTSkXxjpsiIBpFj3R0F8PMJG0tiRn3lpVyVDSLq
CFAq/AywOr4N+gH3UD1Hv1ojdEMNT5sfnc2OewuBBC1+3MiWH2x5TlFb/TuFonp2ziSQGAh3W2cd
vPkzugPadrn/V8ehZcI7Lgj1WjjTRWZmXFj85pmGX4dbqjRes0OKj+EANucFk4U2jOlf4Hf7WRrS
tN7KiEyujtzuuxasTR9pphwkgp5EOlaF6loGdpazC4uPze/m0hCvCy5Ilnc2ctLFt9P4SV+/rVNS
kJa2KFdcG0xQjGKV9Dd676Y59dQrLAsZFcq6YuT4bA0oAb7j2iWzHBphpVYtohkWdV1L7snibfBA
S5ILgfgnZ26OgDbHL74rxLDpE+IvE3uNNIpT/GPAODtqnnHREJi08yCx4KQNFWXFgqmQ99I4cD0Q
atPqv89T1AM9kJFxu68HSQru9w7ZW27w2yyhWhZ8+inHbed6CHevuDiEA+maTb4uUeoPO+4tWNfM
s5GzHJvNMG57Vu+19eOcFFKyxXz4e8tAgkvt2RZ5AWOv65IAIb7lUBX2YAkxZ9NFOc+c9UDDaKyQ
tnBVrsTPDtt+2TNH907FH9zUH2SoK57z59OYTvo4FO67NmrfrWP8qAH8xzUaSdLk9cnltsQKtkfg
W7IM766fdrfUVWdB+3C3vGDk6br45vBFuPyP+Z2aH/tU9be+n8UTX9xqlLXUlXJgrQDXoOQRabZ9
O0QzfgfSpRTs7SEml1BTVtbHo5oRt6JAFVkxbzRXjJIZUAfQNuKePiaTXlRr5+b8JLN07V785u16
St6xxj0I6DatOrcZc7Xu7XahC9Nftlv6pZjRmw7USzz21KVfxZPOqW15dU3sWZhgQ017y8WQZCwC
JaB7VAqf/AV/JuAuGltxWl7gGWPjAUnWi+SZT26OIi4diuebvgnplaEQfky0ihNuYvWApoCtxlkE
We1vyKgxoeqy6amZczm+6xtxMWPUt6AWHkJixur4rXyiOWkZLrx9Cm+AZRWCmIgxXlNzMb/diu7u
CD54Cm2bBTxG3hkcBLzBSEgBsLDiMWDTBAPA0pp0RKuwvs2s0Tu4/PweMvRxLRMKd8XAVin1cIju
WfNKUOojJroJcyqteRdlt64P1ZMTp42o5ndAJG4hDMInSLepON9VKDqbVYSRMdVO5KcCcsXbrSO1
q+d1m9hdS5f7DIqGcK1vcSOJep+zPNGU/dHUSW5uf02YhM7d32s8Z1RYzMJEbD/CmfRFgMI0COtU
6yrHT0mIQQmA/skOdVh18ThYZJgv3WqveaPqptcUKcJl3IXKjTvfKYHlmrhGSOcV3vJ2ythPglG8
OWjcamitWrx/2PiKQtywc3hiZKtQgLIU5aZ68J5LKK3fzBi+qEEBvjJXStAY0fsU/IyrxHbnJ/N8
Lhc8uhXiH6WDeENP/nwLceS5fvXLledW0b34pB01kOZtMMo3jAHKsjNyEgVFnJ+bt1Sx9d89Pfb4
hp0khgSqxgMO2ydEufXvEIP9QXJXRFh6/rDCuEgLNem+459AJgIYnfeIrTwTJjkgUZo6cRQIbrvH
lw1eP2MVD3XYe8H3ugOcBpHfoNVPtOYkiWum1NGZIESVqvKS24lyJOzFLK9NNwO2HfGWYJ5VIwuO
a/Mm1Oh1NhcONIKvEJInaLjREbXN22eb21u0OBI30jN/a/yjGUi9pPmyAeGV76rjsM6FzEE1gDIK
3xYN74SJ73J5lsk0PByNbQhG/jXdIYZuUJTdetHvK321owlH0XZW1xfLyiCfIxHow3hsj8LVwapT
iPS3hbJvv7i7BVxnMhSskKjMWvSwzmGoFCOq9iU9qkr3nGrRw+Q776kvIq7VveFARQ2+4DAjYyMw
JzvdRT5G/jmxEqGj0JDMqemZjM58wNru42dqKI4k0wONrxcmFNI9HxKBZNpaU7+WvVLsYMS39wb8
ESih6aEWobr+I9wNAAYJQjZC3BxMt5ejLgbxJVBbwAJUUUHJIBBxzicFgOW8UOh1Njcs1/HnhSQV
4VrxM1BZ2E69kuozpyc6/u6YhLmXmtzjt4tdobdO41z8lZjA+wCBFVkl5Hb1pQFCwr7SfbMyFyOr
7izl/Xx0HB9c5W3If93hqfmZJZaOWCyIlJjabLCqPXxlCzWv2+olw5fToAykByMFRlTYdiTyIH6L
v0yOBpCycsrMARH1aQxp5pINqT8FRzuFFBgwCCsZGP39cVJD9Bs/6WBJnblI817RYnMTrS7TFv7i
JDlcjW2YizwDGDs3X8l33TA0pUlr97Omc8pg0vdUkcKBknls4PFqZb0ZolN06205rnDIkWOGC9OQ
Iz7YvkZftZqvW+2Bx+3CzAiMkkrasMo/e3BDUSQcBirtHikvk2BB2LSzraIl4AgvfMdjsSDB6ixb
gaiSBU41qUYPUqzy4AuPbyiULQJqeDVU4moRd/pPVoZQrX856pLe9+Sdkv9kBsiu6stCWzTQzfIj
YGo0Y78GKut6dtOYruSonmMZtpxoQSCME4yfIYdtoioraLPGMWELW2k9H3ey6YllCU2/dssDCMR9
QpsYYdDfCmVYLZgAF3pySm2BJWRU5ze+/CAfGaEqR1BcGPKP6SoKJeviu4xSlPMGctvX+lFSXpdF
wCJWoXe4qLxT006I1gLhXnooqe2A40bzJKbMGZkETT+3RE+4mAONQfHD46LOsbMMDt9StzSZyFJT
Kx/N3nMrwSShtN6nc3i5gWjz0gPLXhXz8QOObLBBZkr2uYl2rnr0XZ4HSLE256XOkIa9/RZxFlWs
9MGkqkeF0KQmfqZxx8WLO0TSm65CUPP4v5c/W+cB6UhzQVH/fjyRlvBeghok7tMkZDifERiOSXge
HJWFXb6FPX+8ZavaBPotXPWfOS1sfPjMhHultnWB9GoMw46PHrUocyBCTNl0q9YNQeJf6qqOJrzv
fAhd5FjW/7OuOUJLBvpWCFt/GrS3UiGjKBAmTWOVkKxQRE1ELH3feVvbnucvB1Ui/xVAonWZsvtX
iN35w9CB/IW2J7Nw6c2i88dwsLQ6pQiz9cF6jDvLBua58G1kG3tMZyiPKVgZ55LkwZ7wf/tzMLjb
6U876imFaIgl7jBxwJMqQ52Qwz3JwNOnPRxjq2xmmZuJXnWixbyBL1BvGk1yiq/ej7svI38ezwQr
0zRd/gcKNRe8gdK3d/CMMiLxvnwZzU2nhyYaIoxIkSMvEcxWecipqsUhBNnaqTrYIWa4iPGNrSBs
nFc3NuqreOH/dBGz/RJrXJCDYWWQ8vpYuIvNXuNNif0k9qTcaBy4VpvgveE7JPkdRZl+yRSrE8tZ
nIiRVXOd/N6SgRrtJEOewRa3GlBC1V3sGtoNMy+AYnBhQQ/fR/BI5PAuV7EZpp61sJWZPvtFN1+E
PPG3QCn+P9PCTGTuFYqv1OUf6KSfqL5+sih6UNR0l0inPv2FOqvpEnlCGrib07CTbQfnxweAVZZl
veqTtvPW92mQQj8r0rsNeyZk1PfI+IjfRjY8XQq9SQua++Zavkhdp5LC0RroyI2t9IhLuYV9oQ9A
xQi0XEbh80G4LuThX4ZJkAAydQEH2dsaHf83YthLW5HTw+pha6yiiRC8dETN37zA/grUQOn+XHmw
QtBVbQWpT3OkeoH/utzuQkHV8kOqWYRrrmODTwCYZf+FBqoBd2aGveae4gcZKTrjke92PHMW+Z1w
P6tDdm4wMDvaQ5F6GZn7IWHLvZkea9sJOE5fQAd0w6MKUsxaXbniUhOCEEzgQRIf+ORjrHM3/xPH
15OAT4opdeh6SVWu9fW7DJwPmfZchR7smsI64ITmXxGos9uHCDgVN6Zg3t6I4EM8sCCBlgB7PfMC
174Opns1o+vf6WdIPHHC0ja2HMizOpktLFOPV6U11Q8Ezuu5p7aUx3zv/xZ6w2njqdT4AOszjSsw
RI3e36YE1zwHkRUiLeOesfOOfVJR1NW7FrvN4nL/PscqGz2+vo98nzwJ/KQ6lMjzS2iW4ok6LWbB
tpj83gB9dTq9vsUrLGzdRI+SqLX3tGauHRuWcUqsRlb3gso2gaPEvL567UxbZP152+iToEfcAiem
PvhevTKArw1DNdyifAN9YkEPbTEZLCBb77nJYkkCitdcL9xsfNaBPxUkmCiHZG81/AnkENL8f1gY
HUzmdNB2LeS5Grm1fwHkH/1nfHYyZvVTN2tRMD1htevc8Gl/BZPyTnzT9n4t90lkSLtxAudcWABg
UgX4XFwdiiCZWnxGGjI6QcHk0JpAofqT4DpkKw6HakTEAuwshLL1KaFzTHi9m39iCrpFcURkGXHd
e5OaZg5RO3TpWwyAPFenyGCYDgoi2+TnhYNoZbTydNwI3hMxBw1Ce0KBb1AsZogB282d8oR6lOmR
QM1z/aeg3D9viE7WZKr+bqLtgNLA3R2cwVsiz2eRgk/c2MFUeKbE0G4dxYNMhrq6SEvDMnbxTmON
GykFIgMhvBPbANJxU1kZ5hvN5n+uUt96a2nBLP1iQx5/qr+NsYNBenAzh20aAAAYzmtGhNaXWb7o
v5U7FFLEoSetp2E6/VAwgS7POotdcpBP6+dXN+3TC+SQBtR5UP5Hl3c18nSCc3ppY3/YI3Mh1ki5
WKvbkLn0ypJGcEW57gGboZNyPpxhND6I8w/zNzFDbEWKA22i2R/5uuaI2YsgZn/0ux6LbqPkxoTM
dHB51W12q7wrrKCmr3FJIhN4CfIjhfglbswKnvU7oUQYgWGTykXZh0QilsdR/R6aHrobAUfxRX7f
w5QTZXGoBRJ49LBnrjQOIg6NbvSkAokLeVAk8t7y/7GOX7ecFZtoeu9j0ZqpxbqFClEjZD8fyb0f
HHKIUq7iBaHJH2QzqiMkVe3RynN7A8nF2jzGVr3Y6mWniQDC/edo90eAmeGVi+RU0Y8sB4QVKI5S
l0xdS0gyn42mwGjt2ya/r4biqC/UsZkiVhSNT+JGlN1FL2BVWfNqdkNudzurj/w+rL15EUbEu+XI
uVvRBXf0WNVioLk/rsHxBHyI5jCo7Z7luG+Ysy7euSDIvAJbitCKbBohKNT5hYj/a8ddBhiE/kIE
7ytq9v2OkRM2+TP+XDf7DAVjO7AzLNpfonzxynakkgI55WujfqV5ZlWI+Imxh/umgPS8+0+SHfJH
4w2TZKwWqrtS0fELv5s7Uua21sU7i41Dz9v770Jek52/Kuso0KrfpMT78VcrvwR536fvMSkbGv7M
iZhEGdJXhui5wxro1YbfAEO15kD2vDeT3LusaUwUQVQlqy+i2iYYq2byAnBG63c+YB+KKI/IJ3ru
j1BYyt0Y2xBl/o80VGnr2F9GappcRjpgdtt4l/R7AJxMFU4lFEjZPzQutj7/Y+9qnhlMb1pPKTlD
u4NhmSIgRu9F4FGpx9K7Ho0BXwNRLqDznrAG+E5tRX7utPRNnOq3uyHeU/E3lFadY5THA5e6qPIY
L01P45Y6+c8wE8W+s8f+uURg+rmeqprjDMGjGQnnIb/BlMoeDEvySIqNXifsUwDTs3FSvD76lx19
gOFeMNpYxAmpGXvO7RLPJ5DcuCKU/uqnKfW09PsI71vaegnpQ69vPzLpfUyYu6tWkkQd6qw94K+o
mQv5aymLtjpst1pYJ2lWUqZfpidmSIvz+D64PrV3wfXtR2vKJoBE3hZtovtAn2L86KKdLocIaMsd
R91oeCG0TjiHO+jKpyH1WxUTmCa45opijzFasuR5ENhzD4u2Z7XVtf31NciFBHD8EWBs18KSei3o
bHsfe1QArZ7orIbBqLMOJUm+SXBhf4vo9ZXb8AgMeBf/MRebd+QD2A4PCqRcntAvDaGrhdlWg4+2
47AAs9nurk59nG6ZWzhrYvBTdJ80WEJlkJUT4iJpoCdVQEQnN1Nwb7JaBlnY0XeMdBPF8wwCVOrP
MkonZiG/+q/YAFa/GYfddTGDgSS2RSYJ5LvmESQLImM3rVSasXyOZ27+/fj5X50EHEkVnTyuUI7a
EGEMN29srZ7KQCXSE5NdNzIHdPRYxmIGdTl1EjsllcO+PEgdw7+QHcqEUnMlnYcLmw7wAH7QWCW8
H/iJ5M5JcM7c6ldrgqEGs2kbPWGsoS0qtIShVcfyJSbdQgF0ao8TPxIC1F1lcJjduz75PQcuR5ug
85chZaVgd/mqcfPJvOpgXfUEM3LyYCOjftDFiybpIeY7Uequ8PEJKNLeiRTm114paW7A1aXT91bd
vO2rsvjiWxSzWytPlyBxVzDHzx7ZylXhh+xJutZzWvE1gz2zBCUd5ofeoG+zkUqKveODj//kQPar
TC2aqpbBMb0HxWmca5du3W7AAkmSfoJ/bWAWl401eNyI1urg1dGTJOL0+IpkNwYISJzx7bjTjeHI
QrScZX8qQkB8RqWmEChHwHCxeBKXa+SxoSMeaCZlLshMaqNhuwjsskubAMQANyFJ2LUA3AFvdq9x
nHXfWWabWBMniIIrXUUbkANRuqYX6PihZePOJEDkGd8nLShMCm/3AZIXcxXhOGx3b4zuwfM1njdh
KlMaU49U0SQGkn27ZdieIF6Y4yHb0dOzyB6tlelSFxI8a+6F+uiEIqZ1p2gnIp/hfI9dZ89BNFLb
uQJOOFxVHxSxXvUT0Gv1fndoEQf3TplJFuKxM6gr7qt3c58k4XSD5B5XcK9AWNyc7Cmh54UhLYOS
/HMTRH3fTwr8Wbk6Ga411MTQDrJKD3VY57CRePg351qHOT7arbiTXs/fp+5hORPWMBO55bhb2b7V
k4VK1KzjgtX9RVZajdkj2ThmTwm0HhSavBlp0woN6cAs/p6mQYCpMOUqh6LZJ/Lb3U79e0BVKw1G
+q1X8BcY2OVg53Db0UKDnTy5rauYGLiovKAjV4+8Fd9CDWyg4WEmSVekenCMGQlRPBunrrZMrHZO
NGGocskIhy7I0q/PMVSS9yu2CDnoA6GXRLrazd9RpVAW7sysORNt64zm2vNFFtI7LW4dzX1M5hr2
szJnNFIMXkyJM8RviB/+JHAB0s4nMoDjGdOgaop1E207yxiZ0GBj+8tnXmSSdK1Ue3YBRi9ZyWNL
UK1FNpe0nW8VYXjUJT1ud68Y/anoFdbIpKTRvqUmWHmsv4Ny1zSS2/xP0G0U+1o8RGBQyulMulXM
xrTJkbWgM7Np+GnQEKdF6svJ9U1nhAeSWPmMozE5vuR5swtB+2At426li/CjX99YV7HzJdQKvhgB
Rmm9j+GQCZBsur0/bMKgE/s/b39sc0xDgIVmbbpozEhJ2JNQrN18LgZIBtzzwwDqSuFitK8g1JF1
CGw7id35n0VkHRnDifBHzNPsSyOUisTdWdPY9h+Y92zMOPteVqirVeyvfxhDoObeAGZdstxnVL65
fEtP45MLzGkwkT8cbXNDKeokdslbfUMxiw8umdmf6R1kcqMmlVBijIoDp4v5w97AI/Bqfr9yLwnd
avYgZ+pfSSBQnuri4UUNM4T+Ngb3XdGTqClTv3vVLZebZkgMVbmUsZEAa5frpLTEZ3CMkruZuyry
ocXhraM63eSsPctDFtq/BVFVDrs0zUbBbg8DWKOBle9goh3r18zzNc2oaoJYXGiAtvbULoNC4ToP
C65+xLU08oyqvo/vSjI2gu2meZkf50z4M5BelS6VXyC/vR90q8O7g7DzHZr8xhE+oYh8u/hQsfd8
6CAaB6tztXymtc556OiqBGsP1F3nsMEK0w9vSbH8T6bobaSo9PeMkRkqJJI4kKiTXqwUgOOp5IKf
7QCkA+ItNRPSyu1kfJw3HOjMOGbOG52uxYN+Y5TE3w2DwtYjXhXsp6SvQZ5i6H/JjPFro4i8h8MH
QVbEOeZN5G+YNUiM44r1B5algZGtMPgu73Cu3TNwJDRTcW88xAtHV9H3GFn3osesBeDwvRVB2AJ7
5MCS1ZzPm9Db2qARNEL6wsiiJHNVMuFNkkhYXOtySZn+2Ticjd/9QHX0lywbi+NIXwTS+GvMUVuz
+qK+803x6CWuYv0rc4/70A9QWO0ZvO0rkVIYdbqwoD+AIq3yMu/22LZunnr9PU2AML/zp8+Bmnhm
t6DsncENAQ7nMTGcm/UmVDUCtVuAvh4FpceJgtYSlyde9PGw+Mw1slZyvlG/8lVTBkxB07i2mJIi
tMTZEnU5Pt/KfXcXDw3IAx9eRhDGyCVIaPJ/dXWhzypK77ajN54gGyhTzNJcuXKcG6Tqtm8mXXew
IdJNDI0thdt8TXUTIQW/YEFRZa//HH3+NYs8bxkpZB2DJRw0ahCC/QSen2FMx/B4c40DKlstmSyg
HuEwex7Fu4gsMk9UpFdD+fKj+HQo3lRCdIv24V4K0jcPe65nTEew8DHZdGO6W7LzyPXdVscKITyJ
fr3ftKs/VMZYo5pV0dlHFi7yDPO97IIMXk67/a5cPUcUoq2/auGjmniNXQhRVto8UqerwfbkNlzA
P32sWUnNXtd8CMFx/ESxfgQjt2C6X81Ca24Q3WioWq6Wv4/WVOnlfnggNFneAjCuKLiFU7km4wmj
ScCDQkbymAWRGkfmoVyETenIUXsR9I6SBNFuaBbNemEa0iN7/UnexDQKHwHo3vn8idH6bk0nnCz5
kCEc+kcwXcopXpxd0pnVH2CfUOkQvvEM6nBg8vqZLmPJwi/ipvXwyGBHlqh9Uzut5QEqGyVmfRGu
pNrPY3fCKNcDAX1IjqnCnlhgp2tPr3ybgua2obFkbbPfB19CzcrJ8H1HN6OaIXioYa8mXcSPyEx7
QqfrX+o4CmyPqOe/DVwUhh39u1VzB5RTg7GlVisoEvyBE3BTRbXzzxApoSe+cJqc/r9/CSK37cc4
9rH3Lukvw1pGXStIlQz/5S/lMOIG1Zczl4AGXpl7R9t3JGLx3yhLvTBMi+16ti9KTk9gXto9vV5N
6T+UZ4fe/3aaotO+gu+WHYUfpWSTpiWZ/9Zh4YRlyetreZQKvRKsv1Xin6QQx/xzXIaD88kt+L/G
jxKlCnXfzxfJOsc9yLai3g5m0kHdISXBpGvUxbA20dcK5pLmTmzVqsYwvkajoci08UsV3Xi4UkBG
nBEe1yS3wP5tGCvASpSB7wWPNvwxVvDLThQ1EpFcYnvwytPZOmDh1iBHZR1UzipO302iYkautQiP
MGRreJpVjF32JmYm3T4zL6h/mj8do2qUPZW3K24lNFN3R5FZSuQSFRQHOHXQB17arRSpz+0Tm+HS
bZ0aBfNPZNpkQScg21PaNGfzQkKEfmViHtcA5h0E3pXFqcXwxSpKDyWEdtkt5KdiNbIoPqU++Ibo
XrHWQKX7jRha6NFMWWGjAJFV18hp6PLG3VTnu11R41p7xmr/2OmNnKoc3Jq78SgWMQQE6oacVoD4
VqvAEtHQoyJOH7UIwOlbpw2zWpeyuH9VNbvC+izrzBwiathq2S3xhltPvoZFJiuf1OIRNFEpjdYO
TSzEJWqjvXqWqIHVpoXQ2sRfqRouciAOfIVaZ3OHT98yMjhQtrktxqvnHpnXOJAQL4EjxQ8EJ1ew
kLrOngEBeg+cH4tehT6OzLsdqHjqkWa/tBSt5om8V8ed6AAzbaTXboE+Pin41s36FbGoXuZYYg8Q
IuEyzr6XRbgtI09qePuAuilPI7T/Gs9CEGRvBfxmOp2vmRvetboFeMbhk8BE9IMFKcUpmYFgRpbK
a7d4740D2kB+DIIc4vSMBA69KONc3ZpsbvKqLP01NbWbYuPHXhDhb80L26QU3QrlZy79PCaOhxZV
GoHQVujXAGwKgMFWohOR0n87hoPO90brm5fvbUnR7FQxCsy2kJCe6p80OmFleEOYuu3XiEWPIEya
tVTHKvRyEGO9tnCnBp3Lhm5tElDNNlV8N300phlzI6mvGqD8q2Jluk7Dtg/vzmAa+CGiVFToveT8
js8ZE2D9/1sqro53hhTB6lwx4bm85HNkQMQFLMXWsgXjlSrkmJudsbMs0YXX3rLmprroQTvHQlg8
wlrqLSBSpwQhnMbno+TdES8+2k/F+LO8mGQBRRY0XpCTVbGIKX1XoFu+jZ2ou3ytpqXBXNzlePnQ
PWDgCXebAbEQvZ/VrMFO/a/17q2Ba3gA51MDMbrVA4IMvUdxWSrbEiY5O9566aGp53q9miESBFAR
XMhSUdgKPa/gO/IkwfmN6DMWvx+ClTG2xWH08nSQY4oxlOLUodswgDGDDCsnz29y5jUgaBMZv1Iw
HxlT+MaQoz8YqEwdRal1EYTURVdpXB5t4wSr4aEl83ojENlOUdoCNJJpVB/T2Oh9fGI5DNaYomeP
8t1sXc+ipE/l3gKivYXby0Fdi02WNJnUVM/zNfb48yiUqxUt5q6xhN+cgJOIcn1I8z8U+rSD0V+z
Mzqn4gz8i1ql+ExPIW5Vnk5ZBFgEQT+uCcPTLgjb2/8e18lez7D3S1irWLQUTM4mfLCNY484xEmm
HsWRGGPSEhcsSnAQP/3iSsYUmTWi5nBjNJcI6RUn2QlRW2jxRj/mCVkeCQnBT2KT7ol25olqIyRz
FeQhm2Oc2UkRukVVsGU3tPX2JNX1B64w30AsGv03Trwf1yY5OD5LU188g+fKfJ5aTYxlNGLO2X0o
M7Y9esFpMGAOFFZ8wikPq9nH3ZyOFw5bc3dNLKEvcM5VZpHnJuixeOIcUKGnQxMWPQu3XWpRp/oX
VsetwEXmIcUh/Sq8D8yXuS5jZPLyrZazuI8+mFaN8vnIUD6lZOjO9gO70yEyE3BSn2R/1xXgZiGj
bHPyXSAizpgJYvfuzn7pyvJa3dL5iWi6+QOcg9pinbyHFFnlmYt2frcfLKxIfrvVN4/b57UyV36N
QuSk3zalw3PBYTW0SXHYrDd+Yvh5FEe96mBFSlx2DrayOFrhlwg7Ke1RbAs6jFQcl9Me49Yy6CKl
pHZ3uvzcVsy2xYnGH/KPdBn3iQBYlu+mDqgAk+mVryitMDUoii8e6/1K/0+rsv6Zp371mxG4ZASG
NkMzIARfo1HhBEYljvsCObrZ9pE7lJijCzTYXY2O/opnboSA5FnmuHRNLWI5Bsgx3g4etNjGIhTB
+YvIjZSiXgONPPRqEm8wdmm26mcm4dIeykY8cPCv4olwkpVes5aE2gNk+9kOD6V35u5KJh5KM5Fc
qZtuQqpUH5gUQOs14HU0lze96e/XBZ5bv7jXjviyI92t1rfIEJ2VfJiK65t0fKuWPeUfy38m5yY3
rq5V9iuLR6yj36LD9Sn/CgNvO4stTMWI3JwOfkMPaaN8Dpwl622uk99a3Mz+dtd0QFT/306/LBf9
ezvUoKknoxKSnyHbqKYnXmX7LeHCRnn/ivP6HXCFdhMGXsxhGvAqo0qOu4iI+69Q9FLGf0DgrApx
E3Ng4sSQxQZ36Tw0Jhwa0m9eZQvw9PQ/ZoOpR9AZSnnJRGY+h9U5iOxg9AmO6/v2cycxD1fpjV0p
uWAWwZtNRpEe6laV/UD/OejIetABvu3d6NwXiuOmw2ZoXpD9VPWHsoD0DKwciGrDHMLcamvSe8kY
4SmzfSdBBKlHbtxXoAV4vvSryL6IBLYQ/Z2BlwWohw1MagawRcRZ0JQKqqawqLYGCptT9ciIl/rq
8ziT1xdkna4JROwBt3XE/bru+9+MMUsSX9DJd2JEGp/OMvJRiIzRs0yEObvR16TY9XL0gzPCFbEB
XX8kmxe2pc6ZDgMWX8QBp5NFVozlL6NddADmGm1e3ibPE2y7rM+2Mc8umNl//tDqpRyogzx3vb4l
h6g4LIrTZDXQpzK9AVFXiXKkZwogY27vUU3EM6jU9d8rM+KNWDPmNSYH+BMUYUz3v31gYhYAR/B8
zxL1JZA5xBdnHLD3wiakpwYblfvnRRMyeb2Z2N7aQxtcNBXS1LNJS+ETfjW5yMrB7K2MsWKt+kZR
oqHLatAnZSgo9G8Za+eWnJktVSXtpxWUbXkWlxZGr/jBmU9ZT+wryj8Jg3kdWWIIWLPoctd25Iq7
zeIVEpeEtZhviCXnqLly/bFfgjYhT1Xt7WxsGfvnJRADRAqMozZSZADLaGklVm46wAoJftakbG4R
W54FD3P5t9WcrKQ3lQsRwLQOAJOOGKI9lhYYtKhodUCdt7P/BDO6DblGmUoS3GHocXv5vqcq+/uc
lcXPDf27LoEfiq1fXYob3o4wr3lvXWiCiP+GJ4pO5B+KgcPQeSGLQFykAMKNWi7sDUfJRhZDd+eE
x7mSYBqt91Z+kaGf6+5+T3GBAyawxtsu0Epg+qmIssGQP/sQwGmBOKjywtMQOuX8WDvsFy92M+58
ZPR8KQI4DW+bKdGH6W75s38wW9os6FbeuKSghFQlqN/pqY9QKYrWOrcDSB7nUR0YrYdLKoE5olH3
RAUX/X0bastD7NFMo59yE9vXhYxrmZNnNI4y9lzt9Y/Y5uw3nlB3h4nVVqQ02VkKgRnH+zMZemAp
Tm1qHkg8/FfiDox0JE4Oa0fLbdumurswdYrZBpDaQzbAVjFcvt6q0gs7GhA0QLG3HGSe6xX8Rlk4
WdX/jtDyRen5HPzbW4Ye6XplAtN640+yx6HTxuuN/WPDLPIzmvm3ZMrA8n06Gr7A7nA66lKG5eM+
+AGpq7cX5U2mDSIfOQTCa8ExFIBL+R5EJq+Nz3q0Wn/M5SaLxq5kJJ0Suat5AC1Mk4OuUrifhgE2
BbRflY1GwblQjsW8qtg6wP9UsKJmqmJwMPYh3VtdibhrV6fsB0fSwOwoWOwGOQ25BjIB3pfwx2UC
Ta3Am1jrjQKx0h49AhygBKb7J7ZMbroLxWQxfKGu0p4YRaJ5ueImbStw9Ni1tIk9VUXnp2vtdxBB
zHx8vOvAYZp2KvOlugJDJuuDBIbNqSMZg+UAGO/RyZCM9NCfQwXf+gKYNDNIQT/Tg+WHXayUmUNY
34CSmEOIyVvcRANMTWsyFj81GInqRn9csq342+quEqx8r6IukMRME7nmrMQTSnYxqQAIM8ngnp3P
gEnyZpozQ/fJ1GjnkEZdlfhkiEPobJemLxcU3CivPDD2lUC5d5fNNUgv2mktU2Vwn72X3B/VgbjS
Q4my2MQLROAvkZbludJjbm/WXx6aDeJsM8EfZZS6F5Zj/7l79lxh+buojOJDTdT5YmXVpKdMq8P3
Ap/HUvDvDZBs5rp2eWKhmzORbaeglP93hdrOO1gfymkr0rfgdyIKIGpnWNNBj3Hd+RsI65XKuGO9
4d4oFl+OT/O6QIHgNRNJq0uSxRm3/Sh0SIisU4RhzOFXnlLFlr3dfmYquXTv2xMxPtYkhPc/tuXj
icGbqslwrnw4MTqIyD96pTCWVZOg4w27F1ooTutKyM8BVjwhH03N2uvVw9QUEiwrLwqYhSIXEBaT
NWzGn9uSu21Q6UbCfrwqsncFjlR0cnNKLt6t92AWHR2e0dOOoTvnnAoYX6pCuZe0suoXMcfnyZdp
2TP6sg7jbOUCqPwGG/6Q7r9FLcV0WAE+pcYYOKRCK87OL2PqS8BI7zyxLEj7Rnsvl8usCOsuEcnr
Il4EkwQ0kPVMWekEaRWP4msth2AAeM+qPbFtnaEgTeLd6xKc9E/w33r5BcI4VT5iAKFM+h3VNIvC
HIbdLuPJ2S2Denep3WbfiEgZj0OuP+ZmsBXgOBYu0j3sIxlAG/a70eGUWdNLTta26uiYxqUUbKPt
wb2X4dauxNDv7iAwzuZi9znAWc2aDz4WpVFbQBriKKO/ZJQKPb/B2Ns/sxy1bFbf6FouCLaHtQ1y
lK0/H2XaWPa8p0kRAbSQZv9ARdtFJ3Jl5OzQeBnUn88InhseX/p1j2FsBg2UBlo+sYMuUTPB6Odg
BeMQSddzs5nSL6cNd8hxblqCJCrIJPT8ARsGas4hwTbmB5qZdxPEBfiVoqcQa3NkJM3vJi4NiJVX
Yhrx2mRoRWQ5ifmvFoD0Lb1euZQxru+/5CZpwLcfYYZLz6TVzSsdYfEKRicjaGrMTvq1+CeLoxDG
SDAGM/0zTlH1pTaYiFexlTdJgcQcXKtl7Nh7vO7//zVn2Pf3R8thCU+MNyh2eZjxUmZt4mSpd2qj
y/0mgHWEZKDW++NWlUh3X+Wq0SsBICd3jRmlqoXiUgJyFPr7gfxxL1b4cTvfj3fYae3lD+/8bgag
nOluFJyDG8Vr0JY1OD7BhMi+FKz32p2NDHeHqMYa0tG2iJ9nu/laTAyQrhT0ofzPPZ4HbUzKPdmD
BeemkKUPHoGLOum1sm5LlIMXsFj7VujzJ9oC5FI3nrv0bTvi8GWl9TZUzWdzaCcEHnCr8P6aAo/p
UEPCiTov1pD3uU16VUfibxy26j+OLj785OynJYPzcNYr4SSKjPBuDMwEPwhJ/hEAy+g38jqjtbsv
9cDeJUfRXb/hnN04l9gnc6XJb3E7/M4LPeqdc4SYR+HCJ12/PlMksfBfwy8QBGOvDjHPhLXIOd62
vXxd++aGeuPRlnt22HMumpSJhOp6EyNWaVGHvp+zm7QDNgPrnEZoUsOJblWPeZWB55oqxsELTQfD
2F48bIJ9d+7n7j8mObafzRcgoeLh76OcxD15RfPzfrhLlMxdHhNR8OBDqwnCLi7H3ejkOSWeSjOp
IofFgDc1L0q3wjzdrCPWFQ6eXLqJuu3MV06Vag8uTrAVKJPExGyajy1afDwAVHggh/US7+zJ63xk
XisEzv3WGz2o1l74a9VUzzliCUe2VAD1w316lXlXqWkvM3JQXGgyEBaCEjlLRvvFvn0SnJst1135
iGnJF1CJNDPUBq7ja9hE5sDVGKuOP+xUA1RzNZkPAvq0yN8zXJ0/XZpLadvEv6Jk8fTis9EP8uBl
P0W4eeWzS8rbStQFTh1PBgTABc6AD4ET031LMUJwTx0YdCkYs6Cqipbotoak1NA/00R9RLkAbkvA
XEPDRdzCLge/znLItkM8WbYT3CPCQl4wCnJqUyk6/8x6+x1OStyZdtbgZJddhOLITndB+AzehKhw
WdrNQURT5GyBJOSifIHiVEKZs2BMZD9eWh+VjGi+L8M2CffpC+rmcUWlVviVA65Po0vtN7VPpvZm
XgVb7x78wVB5Y2PeK+jiRe0740DR0nO5BHdQuPaXk1zqKzopsyZdWVdeDkPy+CZBrxAbdaK+PLLr
VkNmBVcE63hGbvbO9j9oXlUJ7tNnaQBhKDleWxWZS3P08S4qwFhOHQtPwUXB0NUZfflQvIJDmz7g
jybOUIGzjScN8Fin7Dx2nj4yLdi4ol1nEYZwOW/boMEoSfrttGyyEqENB6F8mMmZKdbFrq+Fm9iz
VCBCyPSfHUCeE3mVL4a1MY6NM3BZU1v4JVr9V0DdYki0/fcXPfwSj0KowZrA87Kt6JjeYRGu0zdy
OYKooCf4cLTUXwchpBP7MktfDGg2rWgF5df4Z6m2Z6dULbIqTn6QgNjatIirOTMklCrOgihmTTsN
4ZEZ5rq4FYyrhhcskUbSOZTwazKQ1hxBL1Hd6QbgdmqAzLcC9q6WTPTVY00jjzhj21xxXn+YjSln
Fth9ZGXOLwsan2qyf5cJiB8pvDyKEo85sfqJup4mOXiBeQ1rkibIigSINqE93hJQpvhNpxnoc4D+
lzLwq1MVHgVtj4CO1jGH861V3+t2Bb6G3GuBIWDr0JCLr/9GUCXBlu41nKBA61RyJQGXbuKPXlcn
QRS00uwsWXmZ2Jvgkxer4bQ3aK7HRuZxQfZsw2O6PsYOnbSXAQn6KKv6w4cm/DPwFaR5Xzcb9KOU
hHk82DZFcVnvGtQIg1FUCQqr/M5T8ixkQmOR6h+P6YQ++j+odN1PUanPi2At+d+yOpgu7iEsM0OC
DQ81mmi7QciP1stCTIQjW4/ag3IGf0/cWtiX6ty4KDC9KZyGPFGQ1fGrrol/3zakigd9QP5HDiOj
K5Y3HKhKmTJ0/V/xNm23FN4R3Z+YutW67M5hUTkKn19dNdvXlabfO6kjCIyxH/+fG15BA9Z00Z+e
KLHQtQ4S4KpMl3Alq4cwkL1DxwdZRohs4ziGsA4KH7TBH86w9NQeUNksEBfG+QCohq4Tgr1IccNg
iZrr4ZkJk54xzglJu5yoDWDtFqmK+g2SwldQZ+IU/CHwJxXof4TlGyZyRq4KRN5rGU3JRoEozBNj
2aAELC2fg2yqEBIMpenIdB+luUzTvF5+0/362DV1rTbZXjLE9DX0xDqhmcTCtTfijA/ZuQak8ZiG
hgfMh+rydp0C+VYWxkdvZg3Q7KwayLunN+dPQsx98TxpOYbzzUK9O7C5qnm8e+tw49bRu7wnkT2B
2TkhihwH2t/Etju2GYLWp7HJSNTDfEXO0alcy9K7xzsJPlHCq3w1zd8Y8bGsSbGVFpJ4DrrH6b7Z
7tFTDaKgOMsZYwkPUz/8RRj+pZxiaNXis9fJRecqrz573b6b+7JeKKgZW4/icgO9sun3IE3vY2So
0lwN/5ksIZmEzh613Z0WqdblqH8RE5XxZoe7iA5e57YN4Ef/Sse7Uj5OjIzf01La467Nqz8zvuDU
EeUoJNzaWhsJxP8PWd4FTq6HUERQPFRYv5isKRWVLdeJIpN2ZaWT2cX7cMPJH6UTywvuYAljY0c9
NeHT7f2l6fsCXrlnkIaX+5GD39BxuuwYYK9rRroAsQmqJ2VmB7xgnNyWUO84pQp/iQMula0sYARI
ZEtimexC3RsXnhFr7oEyGko9moXA+ntmipuKiVbnEiQhAekSo1lcFWV04073TgqCH5YgO2bU7Avb
NycFzdLxkH0iD0K6PTlqCVIMVVUF/jMaJkhOrisjrPVjPMOzVTdZvgIA/C6lQtW2lU56uUZrumtF
z980kgLUKuxMccB/hxQif/93Vr7shfuZV8cqswey2kYeEvXlaJh3gMw6b5kkc/wdDAFAlGIQ3KLF
ZZ/+9yUXsz4KpOCmKCGJUT837LvoIMQZd55spGLsdF8xo5LaDxjzgQIZZJN/LDPqIrQfvtSmuD95
el0akkAlYBrr2Ru08bECiyNljx8mW5CgNmRJUk8Yn+5aW1P72k8cRFNCv0dx+R7j+YUAUgYuYZlS
UoVAztgujps5HUO0Y7CH4lQJQ8yVWqnBN9DkRhjhQGh3gg977D2Kdm9mBRYKSfsM1mzGKYK3GjYL
vhvcCRS+YhBkOZ3LahD3GpEfYFFFsw+aiQI2EeRWumYSEhQ7YiYnXwInwVeuC6Qt8U8frziX5xvN
QCjGdONJiLu/V9OWhgRPdUpTYw+Oln7AuA3X9bpiwlNQCka5uiAEkB5PytewrIXCFERF10TNADQN
JvVqsKKGnrZyEOM7pLk9yJxBdUCwobboJrJxSrKjJXvFIeR5h+VTBzyvhAaS9WTjaglATNM5uxFC
ZIiqdxv/LAZd79WhAlgRY0IL9CnSdZv6L99IkmyVHIRIVzqjeVVeWm8TYgS1QJaxPyh0n7AdjpzT
hn1ZV09xm3wFavacg0rw55iQD4TkKC00NETJpsrj8R19K2nrdIp5VAasEXU6hvdRLx9KkwgEebXj
TQro9lTZZ3VUNhBoz6sEZLYiql5Z5jWH+57timQslrCbyq1aVL2DohbqLErJ2W9TE6IQDZv/6iJC
br1sUWukBFisiSoP/xEP7amtFCxFkd0BkvRjEW0sffMn3k6Ckh1/Ba0dsR067ERcovE5h1ZiP+kW
TmbSkTa7RXncUQUa9yQ5/jGCYZ0ncsh482WrLl+/uypnEjevFBQLir5eBhyBC2kbsSQSqYiugiOg
AqJeQDycdquzfJUYsWxxOCalFWrjb3X6d0MQWKz1YGWLdpvtSTa6pxXfNPDlObFo4Strmn2y7Lw8
RrN9Lq1RIRtzbvGS9C7Mhx9Z7j4PFDSlnJDkna/JNsFo5XaKn3yi7k4YhEEohmKTRY/nwvIRttf7
m0aeLNI0mRte2nK4n/LczAesxuPgTHIF8G9qStvga2/eN4Ec4KuUoiddDp0gbOvQS8sy0TBE0qMi
rJkovNO9GTla6zfz6e8y7/Xc16kqGqmqkmXncL312AqOy/xogy/mC/ZQtllBG+brl449XzUBtZg0
9FebSQC6ck4Op/uC0wGyP0T/e4FjOahzl4pGdwCT00Jgvbs73AGbYAcLJrUYRhkeIKOs2ZCTvu6c
QHTaHVRFA8LO9YWaAxkUfeunqDXYDo0/x2JwWBpbZZvKFjIMTrT3fBAr84M2W20sXFay/wF/uWOB
CyYRujBgqoXn088jHfJDq44abwVVI+zqfbdGSXY5BhVx1ImLn6sRgBh+jMCqUxT70I+gIu3j+Sia
eNRG2Yp7Q04vlxadeHmIP4uoHE1vqB2b5tfO5UFZULM4tfkMz49mOpAWMWgM9rexRUEvCW1CyMhA
c8JkSr5Km35ypSfZZyJqkxD7Bs8MT5nyuPMRN9SNxi6++ALl+C7MS+KsWhk1aLs6gM5nHf7sscBM
cpetLe0uGwLmDyzmFk+Oc4pjfAoyPqlQwiN8/zAWXCW/lM1/pkSGzKsEgqn839JCUep2Gt6n32J4
JTy4+RG6xhCo6/pu8GlCAh0Uc5JdMHdSMGqOiocHziJCMRjKOdb7VFaANTjq00lkjE3/k7BCzRjq
dDmWjBX/a6+VFk5dyMltD2CGCifIoKwoR/V2BQJCFoJQCv5lqYkkUrf8EzBIWwnINLMvXarPT/08
ieuxDP58x8t4iKxhxZdY3cPZw09r+Wuplj/Rh15hAsHdLt1X67kpKc7RJ/H2h/iPkzoYFM53KM2W
ysfIUk/jfgzxhOrFY92nF/A2knmD/R0iRgdhlAsVMyVYDLBRM2GuU1KRkGCHffR4YG7NYY0GDlUa
gEXnH9QOwUUvjJU1zJu4gQ0qHj2HRzh5/QL25Km0w+BY1hoCUk9q3vg9suAIXml/bTXyted34X0L
XMPBs4TdKFLtVJqiVnklXwc8uEsLstafkk/ir+1YSrrBCD/yMKYlw6Qe/6pOzPKhEN0++mOzUH9u
zh4XKa6w1/zyz42PUAoqflBsM3WUkOhxS5pLUSkgbXtx94rWdMYypwd+79q7+ZB+6+BwWT1b5Gfo
gK09NTfKXycxHZ9h7G0Zqlua7gSVWwp4POHX64mcemgBJJsinnR7AL+nNjFUjdmWJ9vZQQAtEwGq
o1WCr3mzVfiF7OdNdmD2E7E4O7IcUIOYF8Vg9Q1PKj3Tl67h7O0yoZXShgS59cq2xU/XG9kxdlq0
HTUt4ipVO3Eh/jFyADruMfj2MZTSmHMu8CX0ntWJCLLX9O0VgRccLRJWMm4RvuQP0R0P5LS3gWv6
ShatePKYfBVdcwcj0QtIwArcmf64frEVJU2nyN7u6RyGfoXJteacG6SY8HzzGO+gUzjpBzJCM0ED
CoFNFvYVoM/fldXjU97oEzEPkXuM4eKFddgy+/y0AlW2LfoC5/IB4YW6tYLv7FaqKMTGJh2hrJGW
VE/1PoM+yJ9+W73Yn6JPCEECKXYW+EYwLgI4pi/2N2iRxQZP+VfdD2XYbdE0eZuPyt/WjXIneppj
pWPlSzoU9yulG0mtlbHIvqk3OwfhEfPujgIeGzQOcMdkcKti65lAjOwglzoKNotZ5wPAeG7qafh/
AcsQ0m68bGtxMphnHa+y1cHa5lWCZR98YwES1lrW1thk1aF4ws6NM+uUUkYA0vj7S7/IPm+axtKi
MDhHqwvpCFjG9L1f5kmaUDs+eSgUU6qqLiza1Gj7RGtzgxfonXiGblD2tZvSZyZ/3Jems1W/UyVs
z++YA447u3R3fpeZ+xsH/fQJQOha/EtYysWARWuCkrZ61fcvyDbvSlekzt0+jcpwDQugUEU9CXNh
hWRVvd80yJ3gQ2uHe7z1BDk0XHUiPCU+U7E3m4flOQEllADrY0e1LCWc6EYl93aQxQ18qj47lIw4
669r0g+CIpTighPEfOtM5/6mQy3eNJ2pNXU2QlhvNlALCpji+gObR/YVnIquWCpyZetEuygnQzAR
nbw+bOEVPQdwBLKSmWg1mzn9K0tz7rDTP+wTUkIPQLEXs4Vg8vQtJ1txRKmRJMvcqPileAgGlcK6
WPjFZUdD0IH2v/Ld7tCbdxFfWJujOeJP2RR79tWBcR2eTraXLH9GjLtJWuYSMzobec1q4GLhntn7
A9tbuAkjXUrnc08L7dyessLfY8ZlPyDkYIZDcwaBXWa3HHRMpE7k7rqxTP6zwXP676JqvbPhkjQl
lzIAEVvt3j0auwdownvmd28FD0NIzdJUxtAb7kJodEdtv0VjxWyMVr4smpoRlbTJROzZgJuvJ/Ct
J+DwHTps9ebj/UZJFd5/sdUOq9qxr8olsGhWCSo0dNNrcYB7Wqu+UoF9bULflcQnTz/PDydokcLH
O9hKQ7Ph13eg4Cry/WiU17EFod1ljSj1f1C/HGANYL88ILixRl4ex2CCDkWkhTLr2iu2FNPwS2ih
EOoefwwWEEQv6yATNpM5zVBdCnh/FnsVxSt2ZpKzxDdtF8FUWN2bnYYnnV3976Fi6h/NjFGKWWXA
3UHcRj58dZHlaK09D9U3x5z9mboMkQZOwT87nQ4ZTNCjcMtm+IZTNoyIsKT9xEc8wRdMHlXmR4dL
w7u5ynNPgCUDokjzRGbIrSa3GVsKwvQqO+E39fnUjYizYyMnxQzEuEzblgjdTbkVLj2JSVVpjcRO
khzcdwABYVCKyOx/WSyYF/LikLs5FmAxPR4ONZSdgd+cMm8ufX1JwRNeD94tjd3+0B1ULY0KJVah
paivAF596Tu0H+qmoNTo2PVSvjcqjozQVgRN+SZgBDYiOTqufsSupv0qJTdDBljDjzJ0V7goNytO
5c08O9bRbFi6kpRAMYGMyvrktSAUxatQ0HTifA3KhvVOL2yTE0YvpwkpBNJS/PSl6UOYKQQfS4op
voWUge+R8+n2r26DCe1seWl1FuRcnv8RhuC03ICquFrnJOWptnY3YMDa/mXUIukQpydOsEoEVvgM
jDxQeEeTBOWgnYkVqGw+t9t2MtBg0EPJWz7MSzRUO8h19i81E+ppp8JEDSGhQdz/tedhjd2oPdPb
8VLduk2nAhxnmkorSQ2+awtMjGES8YFMg2EDSbDDl8aaV0YWa9bjwNVncu4ax9O4tJ14l2Ltw7PT
XLpaXraRitc8Owdnc1FBbf1nYZTCCTgCr6WdIduyFD6Vg5A01a5nxJJ4LTAkYhAKChD/wqZdwyLI
rJ7FRSIWBYDXcGr2MsChieL5BWZALUcEfsLVcPxv4zhewaV8amjfJvLnEDDEAaU8RE1h87W3Pt/I
2JFq0ekOawTaavmPreLHypXJl0ItVHSfG3f49VQot9MOD57X89cYbq++tlNcrq9prgOuvf0bayUh
Uim/DueC1hXZ4EM95rQa1tNUN522r5dloPn8+XCEj5fCXdlXdsyxYTwAL2oNmmzVMx4UfyKgYmiL
Mb0c0d1WsFyNFl2zn5Btt5eBoSa+NVKp+VlsM7IICy+G5+0M7YUxAcYjv/MOOSLQdCa7IvLgTPL3
H8XEHxXo6WqprB4gKN3dsOhoQnpmts2clqHDADYDCUdht8shIC3ai7clIUGhw17og6NbA48qFoe2
7jjmbU4wPOJagHg7t4vAIcR6QvUeLdOef2v5wCI5HeaV34NXOjV5NkNXj3Lsj60SEnigLpXT1WvS
DOjVK2QB3+Rcm5AlpoAun0/Pclm54htjbappJAoIuRoQAtcWA39OaL7B5xpZ7jF4488PBSzlL1Xe
ebN8Q0OG68tIw8tnjqtPmruQXsv/A768SxG1gNYscnELrzqQzrGIUCA0b2gKk/wbs9mQ5fpeT2j9
GUGaZF98FYviOPkKux9osVv6Di10R/IuMpjBQdax+ZJMK/hOhKEXsiDFqvBrqDTrhDUohNPrak6Y
KtnvOLoktRUEmvL6RrpQb2rzGU30XWJ3zSNxif2gqGx17Vsj0BV9E7L+9oVMOyn4UBMO91Htc6GR
PpwuFRGMn0MUo4cfC5iNO/p1y/il4XAbGKiap5gmOu/0WOWXl5hHvRtQjYNCllTOKWzA9DCvIcls
0QxNHiOvUYLQ4kIsxOceBCq2Ng3ZFEqIQWMpisqsoYAXB1QxpuMHTyWMMr7jtQBwqPj1+9o49/Pj
dM0VZIHDju64t1XtI7CD7hEO3HvaU68G3RBa8avH6XxtJ2d10kVMWxSWop7OwwYSxettDC9pUVqM
V/JNYZ3smC38vaSylVBY55tXHpmZE4fXy177gpfx6+XI2brCk0ZYDU7yHtCLchhq0JhXXDRQL9it
logbJJxvVTumZbgUQndTbpfQzXevfyZgUmxxJGoagXW7A1yen86cgJKDFhTESw6yW9QsKGXgy0GT
poyIDjYstfbEdfmjAoe7NPvmIzmfhY8hvt2meqagdDml0CPNv/2xRlJ9aT3w6/JaGSzRUOF/eieb
IjhT/t9nM4747Zhtaje1A5TqWoqu8ZdMXostAgKXJXc/VI1ZZ5FIlIc0eSyHyejfaaWXcBMcKT4S
VBpp7Cn3S/BeSt2IYGQZHpstoWqAQ11bqFX3OOIqskHm89bUHVvC8+NKh8zxrg/U0HBaYpd/8u5s
cCkqGP3J3Ft89T6htpEK0ob5po3jbxDwtsLNpd7Vp+Pd6BNcrnatHlQCJHOINk9LlvtT1ro4xwaw
E51fFQZuJtC5rlrJSJHZ5FRQ43qVIh1BmrQxa4BYgQDzJyjP8W5WFG0+uIopEkqdjhsL9aj8G9TZ
MDdZN25E9t34tdozy5xlCWZlanpmVW53aPBmFgs12wHdqNwlSLRLrPVcXYNcfM+esVV0TluMHli2
eje0g+TzKaErYliJMWik6kpLOrLD7UaCOOtKHYoA/nEMFZnIwO99OgK3rxXgm1PR1lo6Fm8R9XW3
xFsQm5IA5ad5w051oDQNVS6A1ydSyqIBn8OsNPNO2V2XHmjEqKU2NfUZRV0T6eafipzaXuCTrGEu
YgrCfYukAxihuuSXB3DSRsymbs0D9cUkkshCbhZb0486/zSe+9EASfd/9QYGMA8e+OF/eg9bLQM6
OcFDtM+1tmnQiUaKfsd2NDoZwb+8Biu/OsP4aUmFuIhuVMo/TGaeAZwq4NYFonGeF7/c+LcFjjOq
dDlh8ZjuIwMkKEh1vtmX7Qt3QKdQnfwFMGu1J/7/DaQzbp/M43UrBNu6I6Kx85YTMDBkOhtgarcS
YAssTkl7A6Ts8RdgAazXTl7Hs6QBH+9R48dy7TrJM9IoW8B0cJVL9GzGj1HKaEz2/nxa+scnW1Ep
IS9x4Dx+L62MJX7YYRaQk4KLEo1yVBAHbg2MNkupu+XQqLjcdL/cMdDKn5IiGeCcIuaC6SOUrZgN
QFDv0fL4WuBj22yffUilK7uMrJ6dHS5xr8eTnPfoJnUtpcWx50SpeEXLU+pac9wJUr5/+eTLyO8n
gkj5W1CnOo4w2jZWuuqUjt7qNdy7NjlwRg989xoE0neOgnZsLRqkdt2UtO7DdbyMX+SB+al0l3xm
1z4CCWLOC/HA3XrPpX8JDEIRcWw0Cw1GsbEyylu5DFgjR/KBRz8oUQGmCzf4gu6W/Jak4WlWhKDj
6Eju/1Fv9Fe0O1RCmXc0Xi/pLxy8XivtY+qCL3XF+E9vNuD6PSo70jhG5hpAB4knTb8b7h04QGdt
qxgEPCwNndz7PKwKoKSTMyU6vpvPnsWEMcTRWZNpse0FMmJGFxgw91gVMB4NW/xNNbOPn1cDjeTK
bLjk/be9QDIZ2O2JN2dYVQq4Bnz3F8iLxyyMhyJIzeAnuPRJa02SjTo5pGfsubO/s5aVbQl1HIKo
bQVeH8BnmGstPIKXR54plLZxk8+TF8VhIOSZsEG6Uc94mGpdYX1PsOxcLBQ/4FqnjtwDa9iiZoQt
d8GM5eSc6+bXd0/WRLVbDVjCZ04r2aknstOtRtOC3Se0XEq2mrqgLGvDS507h5IJQafd9lcVP/oN
tBRfvNuRPcWbe5Cbh5/C6gnlqcQ8LQG0E0qQQcjT6ORQsDK3kVTNidnIfbVlWaMvRHjcuP+3+8ew
f/IuJTsrw8if9vzAKi2/m7YIxcQUCnt0IAJ0ozBzYjx2FqKoGVOqXc28zHkktE+WHLnnys1HD1cy
strwxVOJKWcDMbJdob7zVj13izb09TwRC7DH/yZhp6SqbSkLpECgzNUqX55zMFwQ0ts6MloYVIAI
miXz+1mmcNLPAZhX87DAMNj8rH4IkJdxBXB4aPRAyUbvO9QuHXodfSYEKIJ1E/Y5lT2jcdwH1IHZ
lC7dEYAQyfZfxtYGH9mZn1k4qRgMlXM3iVw7dQ/pXy52hEZcTYFzPIx44qsnc6qw4kV6oqIKh6It
MKWMSHkQrtpmWrCeEz+vreAe6eGh8JX+H+cik6bRk3Zh8jBWN0ATzOdI8jpL71fIxSdvQlPsZUM0
8PaG0rJikMkYxHnWMgg2jIqxlPbLWRjE/Mr2ckNsfiaunVNsvmyMCbrpNgww+xCiMPE3kEV2UY/l
U/Cu6BW5yUTb6dKzvA3A2GHDot9Tu+lRodcHSdKZiZtyDXFdppM+VifLyGqn0NHWGGEqwBBv/K9x
YIaDiHOl63/NrtXdyP9jGdNUbccjN6YxWLutGfQSrz6c66e5m3XKxOcXtyTMXiqExRKIqt2/FDS8
MB9Xz71Jr9npx/htyDWr5MAVrvm2y9Gl0R2m4XlhAhd+WXmTJKMdPwB0q3BSD3Qka9FiER65F5A5
jxvKJQdcyTQrwyzIF3EtO49dxe/ci1fBp6SA/a86nl6PJR6qtZSKsCt23xHk/YqWoSS6m+a7sJk5
IJUk//K+xC420jthkZgbwGT9ICHUggkrP5WZKkvmIDzdsLWSHCdRAfhNg5AC3cQ87L5WDAQXdCRD
IFO7rCPsjKFlfzN9IUqfD+tTlNap8hNiV5bEKVP1uPE25+DWln14HAF2qDTkzmv8rqqrY8jPkb98
xy8OAi9vDa5/Qa30pAH8mB9rt/YcERn9PPXRhFLHOwdMLxq1tMXEZNKf86wNQHnOhpjcl7WUjwMB
xRpLg0DZlejleq1m4YqedaQ1vxVJKM2tHPhsMrJGsVwqV1zsBNctsPpxleaJZoE1TAbMRFqx2/Q5
gCNAwE7JK3jDwi4rM4lp8IE96iurUeEuV611YeHOPp/MnrTbgXG8xApt6n9Z3aQrfnayHN2e5QlR
ZftQN0l7g33CrWzdYJ0cfOB19cvkJjFCFK8weFxz47RfeT5wh10IFL92kmlpf53CGL41+jKNHTjf
1a0g28V2zmzHF5YgN8lBUieZZoS+75P3s20kcpE2sVq9Kv2aKnkhkdQjkb50bfGwMmVXTj6Ubp+j
wsEBEjZ8rdzsOtZ75v0fCnNtRFN0VCD2xk1Tf2xczbSMEsQxFq2+IfCfZH+wZjqF8XwvouAz87Zy
gLwW4y9H6FYNFD2GqPBGGHeXxbtvolkyqN41uw+U1zrcCFmwRihbtjKuH057MWJNzU7hBm989UWR
Po3+AvcVlMhtviZDU7Y3FZUymoK6VFxpBipe0k5ix4gmLT2TfueT6bP816kYX6AouEuIUu3HAF4v
qk1g9r2hLZOfNUt0FI0GglSt7Wcn0bVzyOnbOP+Fl81BAPaNYwUADbwN7/97Zt8tzjt3Q4M89H6i
qPlowjLR4ixQ/XMDocrMyzc/8v9e+WulSnb0LBjts7FaJPlrdGl9X6GyMSeh4Gk7Zbn8bOBXqegn
bYLWEcxblECKFeKX4LBKwzM8PYm8TiRBQWx0IR4cn2hYHEnMth/6FsNg8EjyAICTYg8Oq2t9h9FZ
nccuPKdCOUrmLw2c1gFMRacgFOTkdDYyDWDDl9HkmYWwSAER08G7shFkG5AwBU8ZRq1QUzQQ8xX8
6gr/iC9wgZwFE2THaQzVhs2bZBR1sG/Hc9+x9MC4BDS0ylXZq9FfysRd146ydFUntzgScKRY0BGK
3nnGg/pL74Bmgjv13auRrTfOjlaSHa4w5bXtmM+DkXIp3awjdysm15pauzJSdlNWhgICYVgFMhg0
4o+h9ahRR8KAIqv+oG0T6oKOuPEegFEm7J/xYQinb9iK3bI7+E0vcriJcCGEYjGx6sQJjrHqltxf
XuDziikIJ8A7FN5FbzKdFdrB3IRSP/D7K92s9NRgZumfq6cibb+yMl9ADEVxRzBbekVJRF+LfSzJ
ymQlXHfeQS2kx1y2FjGfP9NTnvdqGN8byHEyh8Ogz4ayuwIpA+0e714MDikNo/I4ceQxyUeoD2U9
ak0kua8JBC0/YyyFPnfeN5sLxEtzrSBr2uvpCpmS4ZU0ua4Dd1RKmntYCadpy/Qzn51i3Y9o4VEq
/MgMh+OFERRUvP9aASPFSmZZLhIrreezMrRqaGhEpBitG8YUKEY4BQhVz0qyjd6GNbCB+KdlTR/F
qgkRytddaGsMvsvacdi837d064APpa3aCSDZyItNpTVFPdJhWJyo2vGJl4ejK7uFlsUlFJnoJ0ae
Bdy6RNu7n4A9KQp6ojZk4/qEMi1BFpH8MYsdEkZTE9x6hlYwOaM100mFnX2tMCaaLev+WpTRVbvx
LMPafw2++glolZ2og4I88c2dRB0HYwyMDPye2XQqo/DX8w9lbLqbojozKQcse9jmdhbCKkpggvgP
dsgfBLTFe1o/yUDiBCyrbZy3WSasCvP2jAm4vvNucNprwznXDNpDggkWdjx2m7SBYQxVlfDb2FUc
IEZ0xIubCsF9XuJq0ZL/5p7Kq7CKrp6H5yX9/TMxzeE0AwRCnNXMu/v0sSPYyTNef9QSwJX/Mcdx
JQZXrjhcJ3oanlKMuApegySaU6mVlERMcUWWBx/ubqWibu3XP1/pgxKwo6c+9UXVBL0TMCCe/ri9
0VGn4n4NblXIUgBeBk5pl+211UJFSl1WAi9H4K2Lp7OCAQ1qBsjqpiEJslqo+dtkgxYZwYivz4A2
GrsAxfM59VYMd0qhtpXynJIGViH2ZJoOY1WqL3XWbpjL7gSTQ7ZNzzh5wY4cqCW+q7Ed8LP8eU2D
OGcpomUt7qIa/57RkfPJM6itAY14rM4vf1ET9amdWRRxbM2B5ynE/psdH97b6+eNn32+hUpaBPJ0
WgPV+IxtpVdQVgAVLtMTAOZM17cj22+nw+fgoxBeFCPOwKK3o+Iilg2lT6QMPoagOBcepHsOTtGN
rH9IdV4Qe+oGIV6rpTYITK5gwIbo/lSGRCVFmsuW8LtwD3YpYPw9LSIjBNCAMvz6IW7ZfQ88IMQN
VKicoRufPW0UsuOtywgIc0h9b2h1zmqo0p9fbOgmZUQkjVOXSFI0k8BjYTfU6IsGdbSugv3u7aON
MGbukeFnAhnjhxG4SqZ9eDyAw/EUz/NigkFi0VBMrwzDjeSxBPQZvwOzgxQ291GLSTScjUW2UOOs
JvEQhn89C2u+VIvn+ge+L1WOa3c1icbkjSVzeMDMf/xS5sVjGJ/QBymELi+rkzsXi3C3Ot9nDvPG
KAvC4XFSKg1moOXJyfzc3QuIXETiMx5qPYz4f4G0c1hdvZVeCrWfPobwwP7bOcgkUv7DxOpTc3Td
U/XuQ9zTZUwZaEsDs9XQebhO/GxGZnqYeGFS5ZH73BO2HAFMcz7OjBf3uOsxpOkp9f7fp6Nq1NY+
5PdwUaZ9UJyuabxkdYq5ykivGTNenh9Ir8y4Y116WOBVaIK/JHZChBZNUQODbFjhN70bGPDJbV+P
brwoXet7O0KUSvVG0aM/NXhDVbXyQPAiPVfpoDP++f2riBiCS8xDrZ5n2HNG8f0szEd8Of2ZLoxi
b8WvF2oNTq4qHybapED2/TJoqH0yDCQy6lxelW8YjtOrBtxCC0PHtkAV9et2ggxhD+2S8SIi9hfV
eE2EsLQ0aXPRFzChae1dR0UJr+L0cQy+kCmRGMgwZVKosKssa8ufF7QRfvjm7NbofSTuWCX3yn9q
Q1IvuApeQ26uJOlPY60gx5QN7ca1TZzAqC8rcl9oNv7Do5ll5DQy0G/U6Sa3
`protect end_protected
