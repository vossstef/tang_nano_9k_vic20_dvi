--
--Written by GowinSynthesis
--Product Version "V1.9.8.11 Education"
--Mon Jul 24 21:26:36 2023

--Source file index table:
--file0 "\C:/Gowin/Gowin_V1.9.8.11_Education/IDE/ipcore/DVI_TX/data/dvi_tx_top.v"
--file1 "\C:/Gowin/Gowin_V1.9.8.11_Education/IDE/ipcore/DVI_TX/data/rgb2dvi.vp"
`protect begin_protected
`protect version="2.2"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.2"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2022-10",key_method="rsa"
`protect key_block
uS7CWFVdzwL6ALCacRdHgrkWzFKyQdRBMspesC9U+Ga6l/ZxBRUBRd3a0xNONUQU7hZp8h1YffmB
HB35SJiyg71FPcs5DRMxMGzrrwWMq4+6Mj2vvT8zw8aBHnYlLEJ7WZanrO5wIU9kk+Y2zyGq+xSV
f15/MbcU8dgAbhV+HVvhMfURtv2UUikGWjk2iaVecdvjx7rBoitSEcON6oX3EPtq22KeJFzKXbep
YY6eHbJWPJOWKKU1B2HYt0Vt56WAW+PfxGqyOIBank/Usqf7NUSexzR1DZtKrfn9lLMVNLKGzjcy
PxSuxvCwCi6TVe+hki1fAgpFDtiUHxGSLION1g==

`protect encoding=(enctype="base64", line_length=76, bytes=67248)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cbc"
`protect data_block
huAzxGmg9bwCjUi4c08EvF48KCW2w16K0TkA3L1lSxs5DIAGvLTEcEyR/b+owddQxoNAkyoco497
drIDIEvrUSpYXvBvcal3RjdKJuI1Xw2yXaKy0f4pBE4VZb4RteunzWw0DORmLrlpfS6mmcM89pMj
6YcvPFNU2gSM9NyFvpYBe30/FAyFI06xTBQk34KyecR8Kyju+tsd0mMNJ6CNuZKvWQfKmqjN03UV
LNtaj0p2fceKVuixOwVv/D5i+w8AtNS5T5FbLxLTA539+oqcJg2MvF93CR0wim/sBooKwd0XPR0U
wiN8qrJYur6Jndx7qO3bnQAgszqPE/FjF78NvwzZAGromIDnyfWgZ0Gt2RN9VYIY9V0kKkUFhJb+
BeopDBqLfE7TSd3AQioq3OW9XY+I1dIzEWCcC58dBDVY1Yd7CUGpf2f+erYYeOXvdXhAcQ5VE9Fn
9xxJzteicGRQhIneMK3Q/z3JCuGi8kJcSOoJqXI7O5TE9n6mImfq5WShD0SGzeZ2sQqDzbE9JdQn
uF1HTHsgnYL+2gHvb9xkZ/HHJZ3BMSm8622EmqDym9BVmQTcPDf58saTeFDzfjK3I7kFflMjKJTk
CPSr95XQN/v8mkt6hmrKyNwkfr9PbK+QCUr0bXuBLkVBiRAtNGAfgJryyrWi08lHiSFsH3mwQ582
vKPoYGNLrFB2CpiM6XJVU97US0Gc4NztnyLvcY8r9w4EKGi1ZZyzxh4rj+bNwzbi1TO5tPCO72yo
XcMMl0TLAjpWJ/nw39tQh2RZjfD6HoeEoHt4lAlGBO009+pz/j9GdURtTjYH+MKbTbmdAlsfqHsi
b5oCV2KbrBxb2G035j+AdGpyf5ZiB96uKQu/VEaxbha8RbFBNoKXmDXVrVLjhF5PtOHbrqFEK6sq
w/5oklTTES79ru0kqplXy9juwLCKX+hOr2e15eiHJRycu5TRsamuQSqSsQ2Er0pDRUux1Jl1FyFp
qhBmrfPEySdnX/eQARsm2YCrZnG/aUnsPIXDfIXg5auyFNxOdwnQOuRyv+r1M8am3R7jMbAqRCBZ
x5dQXLVojXNUOPA/+q3KfFDdGKjHrNAFQSSDnmwfydBhCne+VYMJQrc/y1Sf5xzmSUBWQ0TkWTmZ
pAY65Miab3PZ2R0mtzkft6IaZFolfb9wUnu2gUimPe9Fi/BaNcKbbvDUvxJOBIS9yAxtHzd8/qmL
B59KQ85NIp29sJvdP25KHtKB1iE5U9+zLUuJxemmXv4pAoUc7zHi0+TyfN7NjkenPXQtHWPfhay9
+h+p/6YpHA5l7XN/NG01+VDp5h2vMKk/Sgv1lI8mSRsmz4wxsDqgtkBZWd1pJwuytSvptW1oyWEz
mtFTruroSbLxjDBqSWRNgm0UCNTaHb3kdXK/O4mAoPQN5nPvv6hntSw9YLaJsQOmSG7bPUUUksWY
U1CNSKvW24aMQIlFIg1JajcexeC9RgrfjSg7CJ4P5cR6MqRKJjZv4BU1KFyFqus2HiBl3slgt5Vu
+ObZbF9cRRYAg0DZ6zY11toF3I8AQbaSOaNlRgm9FYSGMaJfJKEmJOdLgS/cSBGqEQ4pbI2IC9Pe
LpAoALoMCLXaJ0KDluVqP7PjFfG4gRKXKiXyuaOPAmoEUhozX7us9sdvcmMMEZd2fwdpLu4+x5i8
fB7DRPTG4mGiFqAnd9RVq7aypDxXw0Nw6pJ3EcgMc2lYRQoayuhG0Pb1Mznb2dOzLdr9oZNHVWL2
9OlTlZul0jyFUuQ59zQ0aopPWqk2VJf9x7OOhA9VXHLim8oyjDX0W3cceRLfY9gxeRWXA8AGJxSg
Qpsbi1khWzwD6yAUEjEO6k7ZmcUD3L12wm+y2x0PBNulfBpjHpAWjRf6DfZ8QxWtmz0TAJpWfOlc
gpHINPmNTRvD+Mdz3HOyGhny/chomv/S7fm0ql0baVxT8j1x7yn7yYF6kkdX/kgkfbKNs3O3DFVK
ALL8L33VFnj326QdOMxL7X125MreWA0WdOs8s4u/ItkbUodljexQmQyATIGgD3bn3IfoKx77dzj8
LWcNHx/4T22tGXQ689vD8g+jqvbZRLjLfr1rP/KxaHi3L3D9olB4FtuTGlOlKeJbIUQkqElqlo7e
GpP8bEoyCDnjsawwcPthPusMPaOUrw3wlgTaJjwR7Pvt+wqe2Ccspj+KO3cHrdPDg72nXm17LMa4
9Sr/vB1msmCYD3TaRIptGQq6A9BQV5IYVZ0jGoxJP7EpPQRyYnJnFED+9iVP6UA0KPbMcLcpQqc2
a//Rgdg6THYpLG+upQ1J2Hk64fk/CQxd2Ay+N7/+tmY04Mgd6GFfKUWFb64bZ8UiB28thHHcEIEh
sj9lmMXuXqVsOhANe+RAPbvWCYRNiuMGcoU6UoyX/YDpkoeziNILckjuUL+iw2LT3vzq6Cm9rd/5
sFTaggtrY4U3949lAkjtiJYcfmCq6rp42UmvVJbv0649/VtxgWjRRr1iuIdUcU4lNolF0/+Lp2E5
kXDfwKfgqvkWdGSn6qwPxj+f31MjkbaisI70E6p/AWaxPfGbpgoi9VC6EFWqRf2JyB2u8+p6L/WW
2zmaWvg8MdTuikX0OShc4Wmw34U3WveJSlq5JRxTYZih4947227cHCQ/mzOinYejXQsqMVyJVjfb
vK2uCkyHGjVsR6t/AGWgCX5bEaY/TKZaJ/TnC17+4WJIdiaEUwvZUjpKJHMaBa9wwmvMctwBnycW
qnQFZopq1DDbLyRsCIbJGTOVRsGb8zX/FSDTknD5yXtd2m7o/F1mQl+DPC8gn/8HMDYInuzpboJw
jiJOYYrRM0jcnmNQscklAlJmD/aBjawJkHmZHCyfrOalXXklrP1+KQ+DYjrsjbB6FQIDEo79srJI
yDtQk52Z7/3gMSBCoifuqmx/uSOweDZVZ9faFwfQ76b1juYeYbLnHDwDv1mlCcFD0wtPmNp2cwq6
IKmJ7EAiE+E8crVPiQ/LOe7bRt2y97Xxdn4rf+x6hoyyrQv0A1Odgclw/dmgcybu0MluvfSE19kE
6RkJ0c2bkN/8qJIX/lmbZWXrrNyMygE2qzazBG6rOAP/MwW1rKAceyupiJarlCXmIjJW2Q6YIqGJ
/T+ZeTvuceQFJMdjeTR/3osxQUpU5OI3x/TBSZF3z8NU9puWFlW1UXual0WWxcaSXUFPARdTfSn5
hVcKzngtuZX6RPAINcklC3Q0uXQRf8QWGFybzj23Jtj45Dr4sVcbcqDdD1aE4ZJVhRqovQdvddli
Cm8RkOVngSppRTC0Wv64+GNic9RhcokjYzLpM9kTMi3UGJ9ZAeoRjYFTl67z8DtkX2qnR1UBOt+5
QUZqb9nrNMXmdcg9yD3r7EZAfZV/cdaCPCYxRu8XNZ9tRUqXBFqiiMoWMg/4u73ZVAKnQGqn3Ss+
2pOmjlX2kEj+aiNAlx12U+ZeQC3T9MzjBl1izFclWuczaoJxCDv7G7usHnFA3p3jFKpeU6EuWH60
fI0A3D4N1d7AyWAmXF+z6dOMFrURPgENiXgOxk0jJkhpKwssJU7qZGSMrccpf/u77T2emdy/SNAn
w4LnDacH1MlpRt5VxCWdnjQMx082T6KiKq+Qa9qqt8bO2sL1d2HCUS40XECLzlEGnMZ9hHKUA6yF
amtNTBY12bhHcqqR2GpPUZCP3TdzN5PGIXOWHgBiF/NhGZsEvao15gdLfuywYN1JTmfPjSVCAb2w
GDIV1G5BaUKlzUweZSiVATFvs+dCm5vtYcwGWeXIyImlhbJt+YHyKfsPWkyhOWCjsmmeYzROjnf8
LFP/k07YOWV3WHChKodT9TUIGYwwXVdqtdsl75thODTY6JbVTrj31Zl9gJr+vK7Cc5X7637UQuJX
CoFw50Io0lMU1qAH/Qjvy9c7x8FBiuz6fqG7J0uFUqgaW5nxeQMNRd72DJwRtB27AA5B6A66KpT7
EoM3SdTWbeeForZQuuu9EIYxy9MpYJHmjvSh1JXNfnZwW7HwsE/fVcdQ2dMljr5s2qEOCA6hqF5i
IGFdMbwfrGf6uvo8do9OVbC9XHI9NRiuWof/PNVa8kuQK/0Sg7gXZhx/KWiXRFQzSb503zU3CBE0
/m9sT5luuiWxBKCSyYHvejFKjky4QngDvhk/nR36Crytv+6gcbUTwKzaeuisLFiE31yRxmtkPjeb
NFxLfAWUfUaBaZhNF9pGXb6SacpcN1TmMuw4zUahTpcJKrOGn+BnOdl1rpgZFINHFrmJ56QhgwSr
ItZZLaMc5so/Ganpiwso6cTX8Cbd70SN1zNvqM7wrMWka4syOY+w750XGaOs5pytqVhVthkWKnAa
fWp56DyE7IggEjFev0YKX3aX0p0ZoupQ1gPUu35Epvs03v+ajRS5hSSHwwTIvMCb1t381U4eofkZ
TkIFExVRvB8XCXpV6sUNRzQ1fp2+UvCpz3P7zTXNPLVStcyVEi0L4BJ2TUMAMxENe673V1n9eheC
TXqS6uU2BOhFoncvkzd+kWay7TsYB4mjHKCyIHOXXEE0IsEZ1BWvuCXfyGwSXY1cxUFfttMSv3R/
yOe4FWtN1tlUInLrslFm1D2jcEJU4hmppeSNdw4bZcdHGxWLlZxT23l/+01Eca45H/gTNNoMRWpY
Up0VfCzApWfZoqIKFIJutNV1DHQqEwiXDfAyp6zLOpGlqOjZuBcd9zFzuPatIRqc7OVIJMpo6Ktu
o3Mi1iCM7mov7rKNvA9BIUhDuLIQK9hB4GW2TY5hfZiQlYb8OKDrVmMmzdOwTQ3qQk0fUAcv7Q+m
DWz17xvglXlboiedlstMHlxsOudbahGriR0UzrLaOANnBYOHwotul8R+gLkcUy+dZ3cpt3D3Fq9d
aZD/mmzERqRXh1wYJcaZ1HH5sFHv6SnZ40lw5EKfFHxA66jVyo5tidhsewQvv3Z9CNCCO/zIZCOA
vYh/zCgUedQJMLwmp2j0XciBSrss7D+poeIy6Tx3JdTQ+eE7MiXFmf0oIcHRA2oDUy0KUqiyQzW3
86TiAk2Xa6E5X5lZZAE9ogzJlbZSVXDQYamzWstFCWKwzcF+OgVoxBrRKcxMAPzGKeqWvG7gxhE+
O2ji/fenFGvSJPOrm3+sgNV5OGjzcwu7cHhRPlZLON/SGHz0u2Udhk/HOLSp7muX5iUZbzbNC901
uBKfZMLO2K3XFPBRiIU5PQa26K9wvzos8WgOw8CZYK/y3gI0wl2zhxIHFdiyS6bkmPcKXDGkaguK
aZxGe4E1EhunPcV0ptZOhclHE8gAPiowKyRif+jV2OxmlvFLvmJUuq/GjA9WMYSPd7SZ4a4Z5hDj
BAlMXhVzdlPwMVKvVBh5/UGinGBnqfeW6Tg33Ow2C9cmc6XZ1kKNSDmVl5ekefvG0zMs/jX7U3o3
BCjmZL9lg+NImKUHuLyZKJoLV6TPTUNrLtTnNpg/pYvJxD1EHiLCrPYCRsYBruAPN1OtdJrEBgfv
7Vwc9hfd/lzUZl2X8ZK5dY4Mqcx/foHIKcU9f4O2p9viqKTuiiNc70/QfqOsrzOOWO5zW+/YKDLX
BkBfjTNdmLdhIWtdmbJl/0rP2c5g7x1tfeC5veebfl4134JcpbWaruDz/eDUq2lGuf11GpHlKPOE
zACiLJDz6yrirJlAQGa8x78ALQtnLwyGNCuvNuT/M7BWMN/XKx40eaozShDDZtXJKAq8RKNdx6Vo
CPuYNbSZ704rGPpDD+J6rgXIop7X06IJZF2rFQhJq2w1hfX/3wv7NXOZ20tChwKoiyHAfhDK0pxb
vKoonaZwyKrWvhqMMzOpj8NVQFdKDjszhca7SA0jmj6n1Ha6xDjhKGCmbfGDZ85iezqvqFi3OEs+
GT0YMAdICcE4eqN3J/Azjjlt5Vjy0rp3o3Txv7iNwU59+UFc/S6tabBFyNZlbmhA15EAZ3kZo+Fb
w3C1issn6MJijFyNm+utcgICIdjp/jcoWbjKwQSkk2hJbZ7e05o3TjMR0oAJak1/EFBI8PjPZOAl
SaTCpcPo3v3z2uYN9srbLr0eUR2E4/vXvoJWIc+0AaVgmFch18QtHOiucOZQZyKMRHg3kwWZLYmd
YB3HZKRAbbnFZHbJlRIQY/3WpJsLaWk8Jnj9UQkGBJXrMYV84C54qWkZbUur2wUluyrLR9ebq6KS
N64VM5pwcF5u15Kqte+TwpNzUtYGZEdNWkeJaAEDBnsUs+5LPKJYRF8DxZdAQkJSP6ZGQAn01B2u
eCO9Qiuz+u8geYQOe5Idxx/+NkIhbUvkFkQLB54hE7fJy3m5w6NBNeUlFN+FidYyyKcE3n6ouwpH
Ww1raSqEea3web3MZ/Tn+pS8TFItc7D/V12v2A3aamhWNf8VU/R3Twsooe1AjEQoPKZ7U/+3BiC+
c9YIkNHvZHWGFrNkXuJH7EAOcvJ+Kwv3wwoqpDYxxawrNsMovlhqpuUYpgOEg3E5Bp7z5lp9VyUo
PUiz8pCmZ754bVJaZBA5DIT7FXyu8EUVAawoSOUfaBl7HUhmjsrLv3VJ7JILrWROUvlVRQBGx41N
APoke+BCsvazOewHahKupLVdpoUBgSWkbyAfwQzg57vpcPMzU9QOddpo1qIeJQ5dy+LZKPcrPRU+
i7phlGO/Bd83su8EYKtzgo9KFwNXz6NR3NtRlfpS3XCiR9RvPHmXc09l+jnqg+rJSj+EXzy0ZYaj
dww8qpWlfQlEeGSaIpPfzL6WZNVvUp2K3puB8vzHG/DAG8Wl3zzJhS1z6YUdibz5ICCRRwNGXfNO
MF58eeFkO7lc6ooNIGkbBgAfyUly2sWWQNWdy0I+aZhFWYzf0ND7t3mGRIa5L53g76XeRAL8btwr
QkuVuGojHGM11+/qM89TbiG/XJzOjEgJO7ej9EZtA+5jsULwiBddfwvAEV8E+PrfDweS6qbDAGCn
B02IaD9Dpt18G354F0oX2RSZn0TE2Bm3YqyQFpPsbIsO/2Q8G4m3M6AgFDmMADd9JELSJG3SdhR0
dCiMjTIswTAkhhIi2n8BzOT2OwDFmz2GhzmQLnkkR77wislgcMLo98a4GTCt0LhHsn2BN2hl/kwL
bOET8FvnSIfGSwNCxnD+pK64G209d9FuMJVjwTbyJLaO2/hpOsWqsFLZpZxpuDzgZ2WSrkFDrg16
a5hHaRX1nVj0kEvZQpDY3VD19JN3+2nuidasdxDAqKAAuZ7gokmAcbFi8vVLUl7TPWfAECIi+5kZ
wb/9XTC44IF0YWj3e4siSWS6Yv6PcwAAHMGgdZmTBEZ4bmlugqjeo/0Iz1OYMCWXQPcupuVifw1C
eb910niouNUVwiDD8+eCd86paoYwPmKT5gkDOrT6+p1rbzL4LGYPOCX8WqscNDTtsaTK1XrvRb9B
ZN5yD0P/ziJnMYT+6rQujcLLUlLKg/AkwNvlMVr7Z4r3em3teC6NQN7UzoPOvTxfXRj4VRazRww8
U7ND4MX5E3Wxx7z61yI5/9khcEAQr0rV75jEKdIy+O7OkfFnQjGjTFjgpIDxwbzdOXT2joA9FqUm
Ri+5T4sMhT3B2UxLfTOkGrDyCsJCufRJNLRUz0gxZbN/hyoeQxQutrBCTJM1/1SQX/oiatKL3GvA
Z692x3NIN3tsSYy9tsnQbXiI07kYIOpzloCi69oRPaANh4x1DyCvoQiI/kF+XilNL0k/xrfzBOJi
rEip1XB3Oi1EnPjxYLe8Wlsv4yfJB7ONiXyl/YjggoZ4n35K4yrHFvdwlekaXL/EP87+S23WX4qi
yalDe3GK2QGre5joC9zXv8DNZW9/19lSF0yX9BXgrS/Bj9s9B3vuBaChZC1WaAlBNDQR1LJGUmtr
WUpbPOPxhB/tUe1BKCsf4WpZRyvz3WJ2r1KcHEI/1d4fIAGkl05NAf3czf+01TrBrlV91xCwVsQ9
HHYrfN1Esy+viC/sTfAbvNJJSNKGWE2O0f2g++Qula2CTW+606+zIm7+Fo9LE6eBgNo0HKFRuUx5
BV5NB/kEFxmpQ2OjlbyYeV2xXEHryMGWm7j+2WwW1Lmg7+fseJUICqRkPh4hl1kOIddR8tkGwXTY
bL6qJvrKyrgbG469byF+uXVw9gNIEKNJE5pD8hxABe9expCCy0xj4HkrsCgCl+8jYS6U5fTkhenj
qzOrE06+LZ3HZaEKf6U4IJ3KK0sc9uIFs1xxmQ+kCBaake3TAKzrExv2T/sStVxnHI+5+Fs5Of3z
u1ulysGENjuyzxbErRU3natFVqPXqcYWehyaOIJ5vslURsXcnshBu7rxXX2IyUL8JLQkDsxdoRIt
Unvkl5up40hqOp8oXKaMKpHWQiorg0gJuMMvd2fAJ8Ouw7Q9hDccCJmwYGzAXKoxWYyuRWN/boL5
FAzJHNx0IxyPeeeuRsTG8z9DLZhuCWrhGxTYIgCenqMOl6gFB9WpMsY5bY5r/9R0rKLmBPJWpPWi
tuksri2sUf0h1h8/kFHzbNqzsX15HkW4EGYEYdXJSGsJe68P2jQ/EozBWScZyzd3E2k/1a3M7y9c
og7/aXRVd/A/QuFwIBpBOg702u6N45A/Cw/yijwtotmBzzxwqcT6G/IF/Jqm5eRyND+BMWMHKPhK
B7zXma+COLpZZdiCEDdWDnZnQ+oC6mQmbqAH6EYdgDCnF5KlyIO6Ug6vJiajQ4RYzgd1M7B+TlPR
YBGbikGgoRwrz47hG6JjydAA3tuPiBaljvhGFyr/6FVXZpv8fcFcXFFff8meBmGO/BHA3rgmIdWO
EvYpmq2NXkqhsQ70VWNUYZCkqWxD4NsD0jaIExBxEYc5l5VwJeY5Tq7ib4+ud+z5tbw7RxvQgnID
EUtronXDb4LOwjG6KGKB8ZwWZu9+CUJ579PxA4lw97xvXo4xtdk35GdwxSt8cQnA1qo8gEMtuqS2
2yawePE+OjuEiqxYgmCLJmktlLz4i8w5t5iagt1SKua/Quj9kEqNfeXGGgQHN9ljUySsRGB1RqNL
mn+6RanvkrPwX2tza0jxuLktcBEd8QL3hnb4trMoo/quj3G7RLU8TZLnhT22cjZPdAXehYU799p3
4vzzJ9L1jHoXW4PPQAsF6tuIIRgbz7lA/TebUcogI1col71kyNyK66ZIXA2+gNirLhqf4shZnT/O
k795CH1XS58Rx2ClEZrMbT/imkDSOIzOXgvTG7oI0tWv1UfB7fJYcgZEguqkGaUB69wzrwnQWsNg
yW51LjoX3kMa4JIcDyNt1MTiT756PVAcJUJolnMUtvG7dvzEQHytPGqDi5R5N2bKc/g6lNdJPaHs
iLnueSSD4KLorVgxsJ9wBg8uR1hZ5wWG4iCiOM6z0JUZ9CB2vRE/qgbecYHKmCBwGlJYxDhByOTG
9VqljwCCr0Yd4VEO6YPR3X2TLygvg+o6w2AmBNzN6xc5XCyjggGZ7GbGmOIHp2214lo2j+mYXlSW
RBveMLLH3bKOWD6B770s0wfLyOQFu8Wvy73ic7bndZpeq+LsNSb/UCj5XUkpW2HQca6bQW+HcvKi
51qMztQuoM+vanSOzmT6cbrhZvID1B19TF+/KQtRDqNUCN4TnZRFIPljGjvET8GE4IQZr1DqE4OC
QYCgPYNbS5uF+7ibCtV5wtIQKeYRanY5cH0T8yOb5WbtmzfM47whZ7NEdcfrfFeCkSgS8oVKXnWA
WhA4AHb/MvjRZ7z3pfocaPSAvehQCF8Tcgkz34Qbz30XdPN4urO09l1kGLExeulHW7X9wftw50QF
G/aomv9MMfulZYGO7RKFgR5b3aiiJysNsT/uZCMR2EtF8r50WQzu3Gc6J6CqNuU87b1JoVDM6/fu
n49oSaZ3EkgozTSlXQab7B2GrPVw9Dxzcuk9g6UG1TpQb5ZoLRD7/vGdFt/mB5tzYZYdJtlVw6Ow
F5NvzFzKz3RHJJFZ0CEtJrvtJdQbXrddxil4GEpDLJGuJiF9sOPLssgNZ8bbWSCNBPPWDIufA/Rx
bARUHMQ5q3KnzJNgwyOgI3bJAEDfuywGZJG6uxoBCe0TQuA0zCPk31gYcVncqSDtgw2COeLbwhLQ
F5oY2cp0ioNJb2LMj6sfk5NvLYO/zwratk8XQU83pl3wkOpMxWwG/wMmVJ6oxO4xWpUPil/2wfqo
CXbuyD++T34UA+JEJFIkHuVOpH5QsMDkRSNP6/lpmfL4Vjmlub7ovPdNtt09gZG1N5xulR1ND1hm
TJdTkG7GsbpNSLoZxN/bpNMbQ4xrHbxx+szqla5oEA5Xy6LdwVjEtYPqUoougUN0yYfvBbKgOQXf
K+hVmmMdWkDwLVsbBU8MFw16LuUhnw5hxLy1Gp0D+kAj31wu7i+gvks5szVvmFPLxyy+0BvVU3G4
xiJ1z8ydyiJMxWWAAWEUZffH7WQhkZ1Iqs31//mkaSWX6wf8Gmr6xCuRH0pR0IE5ahHeHSH5DIjU
Z9b2GKyCznMm7QsVDza8Ri44eUga8RlJzeOOOhteksOIDuq11hcYzpdD6dBSRg2AAw0qGwIKOyIP
8axbLXk1FSQlD0AupRvGcIHcxMQSb1CxMDYYOTw9gUF+XmPeHFPTsoFRoNSOLaf69+z/eNBU3OcL
Gi+jQ52kWa+dRtaE1yd9C5rmjelv+NI/tRwmqGJE9B2Ge0WwiltwRegShQ0V9k+in529YgHbVsky
TByCO6cXxH6lbqKU10pdDrCTFBQ3pVDQRymRFpsGruyDgVJ5ECGHUIHW7aOU0nWWmPiD+IjEV+lY
jgJlDMF6W9/ZDB2HIvRd62tbI1hTLUG8pYYEWwi2ZgRhHgb1QyzNFR215akqg2jYIvXQSYI/my+v
njRUg4ZVD5INiAZXjTy70BvlkQ1jjKqgxDs4+ZL1W7noBa6jYV5zI9oIQWh/Ksm2yNuAHX36MomK
btZx1r+pVWkBbmxL3a/EVI0O8Ye05nhNUffIYGAxfApw4Skofk91STTuKDSklTXWwlmNQXQ6xlW+
8r1utWuz+4mwYTzHkdjxmCRnfJqWfPqtSiaJ8Q/VU4xc/jrPaSdOsglaNVi4cVyxTe6cr7xzrRuZ
mayhZliOSsMHHOr0PY0Dv+UUnIOfAkpfcNXaopvWzZGsPO+wN1NkJKfVXt5hT6a4y3d3d8b2Kn6p
ywLw9uFdfGdptWTEFM7dgEeDXfLe7qX77p2wU71JKZKxrJRA25aXrV0AZFXQ6NxmzTt3Lwo9G0U3
hkLvBWO/5JcLSSzpO2jGx4R4Qt9iRo3GoAqy+ZNkDI/GV7s59ixwNl2KeLZJy1AF/bcQgDwPaX+S
I0Lf0M7kRzTNFhJQgtwMnPyfbQIeLvAnBw28+is37WDbivTaLQSylbZFBRUVONgtGrPyjdFf516b
f7oBT71KxG4fVpDyNwptBigJVGkB5KloovdPX2k8eJ6dJM7rCjD2kOZHk/zYaWlzgrOpq4BwP3ls
gwSm0ffoRT4Fly019rMwTwJ9ZdFFuPLtd1ChRYleR+7QneHz9hDsie34EAiJRTs09DNC8YDLFoxW
v222lEQk2FJVtFYdjin8zh0Yg0m/txgHrynb34ME7RQSEE5gLR4Zba35aqJBdxHdBYwXO03HDtOv
UA+dPsXJnjb3xo/Zuwz4mWXi45eaabaUAFJEgTEfVtR9BneGs4IVLbvseZ8MgTi6vkaiQuPvY3SK
bawMIXOndPIWWdgxqdHmHyD7fZlzjRzCOuZn6Uzt8yP0Ml1SHzSAK5A3agLuexCyrViXIqX0+G/R
qO2beb/zftpJYndN4bNbW1bl5VMxQCSEjdvG6THsapskFYnEerdJ3JXlCj+vWdjz1DI9cf2JpP5Q
WxXechVyI5RLEYfAF4DH5i1425lvNppnLNczZ/eEVmHHQwwFrSz7h3a1KTBc27VELurwIrMCj01+
5emeDfaXZ59zxDs9EsY9rwiS+Zji8XJAboDQXc6QVbVPmGuBWFu31z4HfekM2DsCfWT6wX5DihUj
GjlMqtybsp20uq5xMmPKM8NIc0QotRiijxXF/SD888ChDaAU6+lls+1ks4b3Nd7l2/OjU7xqemmb
4QCj6VB5d/aaKIV+FxnFIaaf/PfnUVeb6vbYSGfaY1IIyuZTvPZlzBNxHCwf+J2ACcLPx6BGdZZx
VRdIwh2FVys4w35R6kgvu1DzOXZLm1gkmVNGPobVlWJioxo4YDzXaD4xZDDkJK9qDqy7LNbTXjOu
VdbEalYBxCM/7aAU0wfzNNEdAgeMnY+w1KDp0IfLWeUEta/Gef3MEcoLMcK1h/clVzTh9eQ7qBW2
xhNbhdwnrbpXNCKKkibzOwmBdjIlnj5m6anvlk1COYye8uR1TVxkwU9q2tcMdlYNcvIM3Vuf2DTp
XqMUgbbiXeP6YSGcUnnhI0sQ8mMSOspiwCmu0wkbrSG/6D88EFLDwOPX8bEWhW1MJQWzGmQ5g7Pz
QSWxBrsuGEEz3KjXIxLbIEu6MUbArhwZ6KkI4CNFY8ZlaehQ1SSnNFcOzLvBuEDezdaq+FmzRHZH
oYruhERMvGTYm7gRscqHtwxTLOMiYsH+keag5JDlHCfcJu47SIzlgiyRMthlMy4eAeH9CEAHzfPN
8FcAcco6IaeaEDnK6PaREGeeAcSLMHQ4Fj2bG8Pxq2OZP/9N6Gu+TD+jldFRskEHVAxu+MXUkrjS
WQb1o09l/9mXxmhCB2leNWi+Cl64fxejkxqPWUnzOyqUNkqLzFGCDg4WRiXBdsQ59F/RG7bfVrSC
YGugb4bDVd7U7eOamBZ1aGV5zlB+z+aJtPM/ATehAfCR80GMvjqIjsIpHWI5oB6d3i30+5ad+rwp
ea4sFvQ1pay4kcLKVuJMbj/mQJMcf2H2p/e7TqXD6fE5FBH9QboWJxZ5oki73yAapJtNFiMtmaOX
MSKCvLWIaTurEkEv0A6A5qaJxMe9w5Pcf0ii9EwUl2YMvNrGsuh/q+jk2kI336FSP9X1nC1xak1w
0835YTtxMkQxT7hmYbXt2basr1u2YSNWxuugR9OUrura6IlG29EUancZtwfAwdo0+ti+qcF2QEnX
RyFSHgctmkpAGDo/u9H1d0tD6oZpPRNbJ9IoypxN5EPsc4hHDV1WNo164/adc6dBKDSvL9oBYE5H
DX0QYhtFIya8gE9NmuCVhCC7XFltfByeLTXpWwsSX4wC6mrcUsG7HJQAFgyWow1HoaO9RbkqNm8I
jBphQBseY/ExdGNXbMtMmeytFu1vLMKFV66t56SUvt5QfntDdDQXdxNf0fTWYRkrH8Mm7jSc6b13
as+HGX/QI62EEO262Cjb+YxIthDIDQ6sltCzkb0sZWSntPCDosDN0/eb7cEAB1gcXNAMA0mc65I1
uvHNTRCCs/7bWQs6Oa1JLv0GKBAMQQpa1vT2EC1F1GaZ5YihGFeA5yG40CrTytNq6xQAkQ48jQ5H
X268ShOoUeNVFJLq59mMCi2wbpV75kmBizky5/Zyjwu2A3TKfyyef+l4almDNQqbyulcVccdQF3G
47CnvEz24v7H+iVJANMFH/P8kSAL9pnNkp4Wf2F2m2+Vzt25yGAlnBcHbOGf0tutKx3BcXE0V0GQ
3yyuGN0KxDTBosflFS2GUm5/+clK+rsfYhQKusJJCyRzGrpg6sncR6WGKuFK+uXb9dKRZDr6bTLW
AOoDdeWtNob9U6R+Fxq7t5fBSi6DY6VP0Yv5ScHIImAdPQOKJ6/wrcLV2gNIsDeKJMFm2SfIiEuo
1xLgulm7c/RTAjl2Hkc8hivuzRZz5e0A/ZmPcJHvqcD/wYc3nQ08AHjQBCoS4tHGRVG0crGPAXG8
XoInRPNNB3HXC04ZSVtzq12gU6Uh7kPBM/fDdK74Zo7KcMxuPNWr65ETUMtYnN0xN2hDbT8IL0eY
Mvmeb1VXUY5OgV4O1DonCEDPRj9R9f2oENVFPqCUaNS4MDM3aaJnEO9qMQ849ubcifeWe+czfDQJ
R9bzUYkYIrqcDIq2XCmgX+1H6aeSTwmzo5IX+wfHOnQUogjZXHGcRR6pJWz0Vzy90Ds/bi1ZGcir
usJL0p2aDdGtCq97r4xnE8jVi1+vul+lFx2Ouo/ppCzgCiP4MuJfB1W50keHtLNgggRyiYKXvok+
J5fN79Bd0Badi9umpQMlNfkxEcb7jTrQydvovfaiMkkqN/xKNizVE71CiIIPgUymuxSsh767tAVe
S9LdqiyZh4wf2Ug8iRcsyqyNOdXYZZAGOw/Hof6Ix38n2xbbnyAbdHXu2GxfgwbZ4UBRoBje3sBv
egBMFj0yJwwtuFIIpLt08dg98cT/T/u7Bqk+4rGVOTIXQiHjopxAgy1BK1uR71CHo/CxQm0I3GaU
qhNFWExvEtZknGzw4Xe1QlUlzO3DFpk/pn+RtliBSDXoEfZigJ8WxaJwxD2oiceOuLFHr2mTr+Vv
Pp8Uge7JUj0ERWPi04MPxD6S5bBDcmgBZAvJ5hoCe6R9C1m6hzbaNqcd0gNuKgjswC6tayXjP1hI
kxfZdcS+y7CURqzoUervP1gR3ZcDENhFslM/VK7LOpsSokxL9gYG8lu4PFEuhZLwU3qoacGPPD8y
c0Xk4cqzuzeC3zu2IQwadzRSCiprVK4EJwY0wSEexIsxRLxRgy36hzGtNgwPX0lJnyn/0c0Q/QS8
eHr9I8bhEv/7tqTYa/nr5vlmXdcZQtBN3iw9Xva6qGpN0E9pZJaC8Ai8yuXytiz4Jj4CJknirIUv
x5ih0jWw1O9ioVWGL2/vZyQZc7gxq9ADyP+36GBiGf07rKofWs62kTOCnnwFdR2lnIjTny+hm3yE
gX6t14FxVtFTdXQXwYl6exaKSIs8gcrgHPGnmcbXB8UV6sSa9bk3ER/+hA0hS6/4XBzDNYBvIgf0
HTNS1Ph85VHVOPrkIrntVnvIwNEdhSRhkKTM+QQhwN6ifeORtXjZ5B1zYoZc8YjAxoJx7wNGdOSt
uyI6cOr/joxUqS34knIe6AYjKo3VVs4BhaE9zp760TscJIY8tBgJm3UmfCGWiga/U/xPXpo9IYdF
QgcI5egtW5czyYnBBXfKlOpY2t+K28ctMifTATTnCI94M8IR7cJCKfTQXHeRzYNO6q6cG/Vd5IrK
uD5qwzyR4++m6UhcBm7ko8u4SSnikN3HRpXVpwCrmRxh6tQSEOW2g2LByGzQD/KVAwd2VbUIuIpt
i810IUgjjJPpx70Cv6xuYw8Zn5rE1bzUHU7Lvap8t0XQws5HM8KSSBUIzNH7OY2OPl2HwfoQYWzl
8Qw3SqIya/LlgzP9/g+8WMqs3BZnBSo6YdikKMP8LW4OFE06xr+DH9laTqEG4y7+uv3W7jGnK06v
Ug1iBOhiEaEc3W/8ZzaIBX3gDqK19OOkoZ2LcAHzVpbymnjxft23TW4BC7EPTRD0nUW0qvOwxpLo
vY1TbAT3AJW8/EhjM0oOhGEhKBmd/36y8S8mSoblUiwVINu4xRzw18H1EcTxMrlwkR65ZNrk2Ong
BjOq2jX4jnmz2u+M1aFWM/O2FV0aG37+2Cf1oUe1dqM5b6iPw3NxfWzs3X9biAJzbov5+mBhV+xV
+4Bmdm2iOp283BfmUvRHU2SLp+nkkrAGFSkMiNLeHdvGj3kZYs2M/6NvgJwTcHtjJxy9+iZ8RtYF
qfNcsE3U/7pD0lxHuaTpliBW0sv9gGnirJrcB59pOhlP8ON92nrSE03tJiSC0yv/0kRaxg6JfJM7
wp4ioGkV1Qv1gg2SGKG8kbQ/YNs1i8mfBjRQjsaMGOYhoLAYhNCtwbCEmH8zRv4R8e6KenBn+HJ3
EHk6abgIvamHgltKYyswxPNEacwTOiVKGu8dRdfuyY5/Lmg+7vmkK1rUFIwZStHVYP+2Sq4C9Bcf
S/03M4MLa8lIWB9o+EoQ1fhvKhRB/bsP4I03un4A9EqI03TU7wIrOUa80BO7pjsuU3iMbh9OHXjm
n6/s/2rGa4N9fU42R87W1vz733xiQks1odGpcJTy2C0qE5KAd0Oe2bbypCdufFRh0dEDZDmXVNFM
U31Gz7HMePpG7sFKHG1IpsrPEb5I5MhRqGvyd75iV90hbVmmDKVicaAGY5X18ZvVqQt6M8TyuVNX
kmqT5znxs8snKOkOPcwsmfDbCb97P6ZtZp3dUVE/Wxj2VJAcpL7h/Ch0RLCUD1kdHXNJsDz+S/Dw
hPMbThAf4Osw9Wd6cK0D5/y/gj8+rmIyUVQTZiPtsYvHmIKyWbu6yXgnsG0umGLP56jr2lSk0CT7
YKM+nW4VIlvqq8zUU1tzjSxhhKhNnvUByH/N/BLwhBY1/TXpY0ioVEuQnOT6iWdnEP/eold/v+fY
ChIBEGNJknjLaXn3/QSEj4GRcdSnum87dfTYgnFCrXcMf6SDUXWdKYMb7zYlpNnep2ALzcloHXUR
Lxgn8FXo6d5OlpC/S2C+2gH8xrIE79+NfJ0+KB+iuiF9+mTLW0uNgsodGJ1UPsaPhtlgV9eKfroD
wpoyUiMVteXJba4aPOi3WYEc/ogTNx2wQzTFft1IjZOEJk8+DLxbcKJMNp6+EI75Pg27mhrAMEgk
y4vSJCbw6ROXCvnZc25cPoDCJAE83O4RIXMZqXJm1XV7eYS/rDkhABgfwOaFnXqojnCy5g77EfjT
uCTO/fAsyGuYyM9HOs3VrHNSVf/bWC6uRcfT8dKDMTqUTG7rgCp0yxq8Y7rvhmbuZVEu6SWhBnDH
VAUUqZ6mPZd6bYsF6I7ePnixuWgTBq1Fsb3CKYKIBNy58OUFXhaeucmOUkQwiNQkgKP45v4zQJ4A
Z/BnFd8wkew93zgvrJGjqnxyoZVx8RBgBOVCPn6fI28vml8nt/yvLuNSqkwSnoUU+FUXNtKU5ZYj
ESGUgHkohSqR1gXF1gkEgavA4/qUm7FC6VtGXXVIRt3KGsc3Fe78b7nvE53dbQQmZ9LOIuvJ1v0/
amaS8R9EZ109YFfxPQRgewkytE2uml/3yFxWXPl6Br9rN+L5O3pIcayVcSaJfG5UeDOYd8tAUhKB
ygRjpD8XSsd2PbMX1q7EteZJszXFqcFFkzQcDBVDbnREVS97ynkA2pneT/YKf3sT0Tx/0DSX73OA
S/xQOjAyXQcqGogaacb3NvZNJdWPloGoaBGSdnvGM1K3r2R7EWRw0UlqWd3b1tuQPKP2sQt2TOAA
AgGkeEQeDN/XyvNbFcYislac3ARTA45CLu6SogeEtLUK+qlyjV93PFUpx4Dbx2S7n3qbk7mEgFHX
PLpf9OHZZ+I+re3ypxgahE8kFE8aFCg1rVrY7bB5zki4TyRpIoWpCE08wcq5RW9GNa/IeB0FElV0
oE6v1GP01UOmpxG+RYdTkdiLCMet8ivWzEhXn+72L+mzzUJzyjXAW8EFyKX2ZV1Gd+ZULi+FSANb
C6TnbKRxiVdTUTRHDVTuQmMhJCaFaHwqcg/Xj1RPkIviL7kJRLHdLYOdWLqgNGaoVOUn5maVpOFK
BMw+FiTsX6evKal6zlQrEuU1Pni0UaktqXQiZ1M9IvUy0owPV/iXmz0FxZHYe7H/RRHyRAOX9qT0
EQTUQ/tfyA7f3AolqUb1q3HK/ZKnVxE61j3mIb2/IO3tkckGhd0IwHkRR+CIzWcdkx+fTAAu1ja8
wRYqr9CuybFWTCo0qRWE6jkiPRrlAcG6y9EROROCb1w5zVxjAQ/feXeFmW9SZv3HRwdcdwRawHcQ
ME/usNt/HGDpLV9eKI8uQ+/GZWocN0pqk3+B/OGEvlzNcCr1yz1v2Ok/mnCpCWYIlx5X7qXtPz4v
oyVr4bh2j8Z/6XRG0DZ4jhQIPS7/pOxePi76o25ZzyDkDGFvn6cLmZ7H7ys3cnI0NRarzbEBOGW3
hlUPtykT6YQkyQFsuXFsREjq2m3WB2YmZq5t7YeBRTm7FVUgFdjSufJoiUSpCfNoE3S8quBN+X1/
5bHslQEim496beTLCP0XaqXJ8q7SLAfzzU7tlBdwNMMqiYFLPfk9yyUFnxTpdY+Q1snaj1julovU
KaOZwW+VK0pDPNjh2HQTK1uIcpk9LdrsiOYO0dLCkjVuw4S77rAv4qglHsSRJwqekLuNzw1z+Z/s
3sqiGSJSxfceQ1ORDvtaVV99LdruqLwVksonFjEI+UbnigQ4EyfIjGNdG6dcCrI7rAsDFMGcfpK+
Lle4gnQuHM0S6B65jSXcqIgLftDFECstSAyjjVPiStT97xTpkBpYsBI74d4YeMTZDrJm6dXlVX7o
3SYBARXgY3SYG2sc4XHUntVHMOse0RdpvryA98pEoul66xImK2ZLoC5hUnoZmvXP2SWxpfZCVMd3
7mBP2+MnRGjbUaLsHnVQp6R9twCpWOxeP+v9N4DaC8C1JbT1RLS5+59wnyjBRXLOpB7epTV5ftpw
wrpFd7yrGHB2PQljZUzjNNMUndBrB8J2t/2FtgW9u0wPPuuR7nnlIzsevd5GXjKIi4brFwcZneMr
ieEq96bWZQBF89XPOL7CnZj6VjCDQysTULS9ZL3eWLu8Vnunh8+ywE9PaDzMaS2rYH/0F8GN1e1N
62F6FFYosc/R+tjrJtMKCADhIxAk6WZ5vQvPzUDWj3Lkmvpv5O4tqbwGW1sNcO+3OSfQrZwZZw68
KntrVbObozJR2Wb3zhr5Wow3iGHY82E1zWTD/CkN6UyfMfDenc7lvc1MXQk0jTIRxCwcGbxA24kY
7JBG66jzP6g3IVrczV1G6NHBk42B8fWBbyV/2LxKyWgA99Y0NPR0aCQ9goqq0bslFJ4BK8PV1n8q
aVriSJw8mBAB8mzkLQQ87048j6XYF4pUz4wGvri8LqvEJcTdS8qYIFI5FpanGKX8QZ6eXDlkJPhU
GA1JTDN6+ZK6StP0a1SdPLIkzDzqyfjH5r3RgyUpIpu+m/dS6humijJBDawuX2tfsHHAhUk+0Ly6
lEoS945kkbGcCKAHgsqU26qnsISYuW1PS0G/rm/Y54Av3IctQCVPt0d2K4oGNpT6QEVgtSqDvclv
Qo57XA16T899GZ+ov+NmtY8jj54mUPwJ11jL3pTPgAdEHKbTdfKsRNgp81wNvHfUcxbfoiYDmrBj
AWfdshkBHnqfgScX4eKYOipCuAzgP/G+p2VTw2mwC6oVY+5miZWenr56YanMNOGUtArrlfo+oF23
b8jn+r2KS8BMe5ZmF23hwpFjKHBhryMhhetL6ABnrjWCQerR+PyU/L9YV0k/Q82bg+loLuslV6u5
aDpnsQuQJYQkfGMaRHWj8f5FeXkTBw78+x1k+w/ko6edOYK+3UGttxgDgOV5RcFbYdfdpuRWg0yK
B0rOUB/ZsEy2eB+xJmZxbzl4x8+GZE5KidYmsPKvJ4Mj7DRdKw4UIZ0hDLFQEJlcMKh8hCzpbi85
i76j/8KvKIGj0fX3ZbJdkPCRCd7X93BFXvpnk0T/ZxqfbBzOoxohdeXnO1lM0/5JOz8gxIjfPXvB
j/Wwxt1sfoEe00V0hxXwZT5wxeizJVjWO68MZoBXxEzwWsXi7xWH6TltG6Fhs7HevuzrNdo9L/TG
aFhqUGC2rrN+fFljbZ0RfhDjszUjAWJUULR+hnjDdegZX/wy0x7cE7wqS+0ZBlaEoEgGL8sZqpZk
l+0/HJNYhcg7mjSGUdbE7qF9qyGxUAUeZVgCqWSmXHjdS3XEMSfvf/2nH3vG04PLtqkvJOfpJxa+
ZEI1lM+aREaliQ4zqggi6IdMQAuH/zyKe2kQpPVOjzZCuFT/X/eMEK0upEzQHtfdwrlBmQ1Oyz6f
DOdJaKaNroECnA1d8AHYjc2IPNzAdfyhQZFLQ4icQMp2fP8TYTVSd+SWfQOCikEClSa+5ILECjiP
ADkPjXogsB5IjlvZF5Wb5zvTDhUs4ZVZ79vFFduQlwTKWaq/fsCed+z6ICfPLNO7hQqIdtnNmD2e
p61moFwtAQzI8ECvsw1JyskTIFN6nLYWaobi4H/AE2F0WnHShFJVWf4gr5sdGPd3uE5UQkdzCUoq
RnKA+y3LrJuGpGm5XySrjGUQpzSqQi2hpLcoDZ3MQxsDIE8CW5BhkkJgQpJczLP4J0n84ESVHkRx
w/LbH6C83qotnUUXMbE2CGC2hAK4vwb1YQqs6ugdXvxycUAFV7TPgW+7q9hMey/J9OBf20i54Acp
ZZaEgxvaZ9aImCxWleKQ2wyo2O0RdEZNcpLmqvoWeprv7JOplvepaFkUkMmpy3oB0rqmcHZD+HFq
FQu9T103bFPivbznIilPEmDoAWp3X4LlZRCu8+YJ3WmFYnK7krWRRzXMkmWS5j+ydYgajAo/+Tyj
JmEfdm6yrqBuct3XrMoYxJMGbjGBoi4bZ8hjWK/d6P/3f8f/bmb9P9U/A9De0DKvtrLoGPGJSlUP
Rrm1nC3C/U/8jxMDSkHCeAbgZ8muBKJlKHISqr3XyrDcZQfCMvRbcAnz+WcicgG9yldwObKkHuDd
QcrhnozEOY8au4+gUMqIJiUcQp7bS4CBXeRGMaswwjKkAYhSywlFFFAazB0MaDCCCsVCAMiNtYwe
LZ0ZCnSrQ9kplFdHADm/af/mP24MCfOjuXK75J7s97mnEnK8/bopkwp2xrZohgJl/wglDwadh1My
R6CQfPRy2JAHaSt+HXjZkfjjcWUHiEduaN0DnF1qtCF8Tv41HVfZbf4tLxpK1ewqypoAtfT7DbYZ
qSZUSsrgXMBWTpRYb/2eVcLS5bJ503If6W93CbUB+cEHYsTSuYyS41CTg7wAwzsn5GlzY5/CNK6f
GqkECHlR1jHiZqQxOHhEneleyBDZF+Q1MlbiCpmrDRSLtIZGgVjfc+0ZDP8Xpj4VNXoB7XHzHcYm
E3cpdQMwum6Ah2TOZgiA/L5fIa4wLB91Yo+ovZrJSb/mG18CPnHcDBci/4XZ5+MoiqTIMyBrZpyM
j9YurqAy+68rfu0zObdaqKMcPTiTwkJ2IincpSoAFIQLWM/R69Rn/A15hiEBq+Idgf5qIsYgUZRY
W79bfcT8kpoPuiQ9tIchSB45nznXFzLRrcfFjGyotJoRImYGsUSKAGQ3b+74FJx5sGporyEL4qCS
nqewoFYhJB0hVoQzGJVAx7Tfv09AW1NWkN6u55IwFgO9S/Oh09wUB3oDJgPC4G6wDY7LUSw6LcCC
9INOXYTH3OS6iPD45HxG7ug6pbxMKVUV5V/9yI4NL+H7MP5vnVhKlEJhJqmYY1brdXUHUsNdAK15
u5ePAK54eI8IwwLMbazKqZvfTuiSO5Fz4cDW3QDvMAuCtlhdizeiOwOZ5T0IMPXugONpYB93K0Uf
zi1MAUFFUo2fDgyy+8QUA04asuoga+gBpkIPK88oiqyb06w2RIyMWBrxazmzzvdjQ/+n4b0oKO3t
wEGcFZGhIBqTJmu9OcJmPtHqKqkWErCGdjVhZotj6RmAHFGtpumB2wlBvotLLN+OTEE1z/e5BJSR
0JLNSCBAqeGcS21cJLGM5R0I2HrjTRkIzvB5RMvv5yW3DL8D88Dzw8Dle1gUP8zmgNYzW2NJo4bT
/ph438gAbr5f9KtB8TVk3VbEjUSAPgqHcbjuYdJNt612y8ZWFVwaGrkJWuIPR4bOMWRDKLl+zrhT
QNGEqqcGc0fj/JYif6jSfnOi9vWIY2VO9LcIcZwofHMa+prtA69U/h1ZZU9O5Sd8tZUKT2tPimfM
fAJrrh/eOY4gnhXAz2EFQjiSQ4Ocm8L3LuxTCiQm+oISFHmM8JP3vxutxA+axGVV29dU7LeK5zlE
ZEgRNrGlUPE9srSoggxiMMhHym/WS3/RVtudO6BbTQbj95veVwwkUrV4oLui+mQvhqUUVtoixmPE
UjUI16lnqIuNcNF/CKw9d1kKi4+QAzE3wfeZjWwd2D5meHn7DtyG5MMn1/HDvcs00eRvaLRstJQd
0pb7x6LhPDyrx0MZXCg/NYdME5OATA/NgWXG2zWQ2g/XYkUBp5AeOyMVg1L1+gGzxBd/7FXNwh3o
kHUBsTNblpOMn+IXXrKd1AukPgXLgObgDtCrZEgKpJaE3fUJ3Zf3YwikaP8X9TjjbFVBptfncZew
gBPL38rjBX1pIfOPgHnCjJCe+/5CF5DdKO7aPIEnVz1tj6Jamkaj7H91KL0MEB7ZanZy8HqhhLFA
LDenTVvYhRXiLXkb57ScH3nsvznPNFH33G7x3SxMKk/tPMIRd1XWD423mPEhTqc+yEuQATjR1lfy
buYQC2XFnJ5e4o9N6G+lpO1mtIRbz3XqzDBVrqoYJQSHSMvtQa6ym5riDOirC6o7trtWy6Ukrl/w
n4ei/jrtF4h6c//5jPyGfzQz6hgT81pyMg4Gq1KqgwCdmb7zdIWSodiBPK0CP8Hr5HJCErGhPZvg
r0mOmz2aqMlHS1MmIhpVKlt7YANJEvlP7GD2llIb4D+8mvlcteOPsrwJQvBim5SMWINiDLj9Pc+v
QsiVOD/6afbkfgOkzLM5UswCLYZRddbr04c9UeSZGpcowxSSn4E0HXcHX6HIGgt7L1Jc5j8EiGcz
RvOZ999X1kg38ORcJMaeY7MMlznliLZUI3MVqLCxDGtGRdZ+n6DV/EAVsJ1udRy6UElt2I0MWkqK
97ZR0sJFCpeXHPTmLhrLbjIX7crwoUD81iWEg18tyQyeZIcmUZEk0bS9hHTclw9YEEpjsE/pJUGG
MHO50T3nfYtFeTXdf+nYei9hz0e62/Kv1Cnp+1Gaf+YviWDwzsUsADpsVgSAkszGYDwkh5nnRUXp
m1kXfKlmq3f7MeUlRENdz8LOzTT2FztIYblGJZHuzQfZKuDTQTRWrCPIIKFI6zfs0HaB87+XzCME
kdXmSnaaan8LBy/M0kIA54kZklnyQ0K54c2r8M+lEqfsdpKA1nQlxw5ktI32ahx/nOGUNcww/1+o
RuJ10WFSw739o4zmNbu8c4RMDB9lORx20zGhDhdIFuBt5XuiTLPa2smnQLn7RaNnuFUe1oiM5j8Z
JXRSm9fDchjMiXPkOfN1eJYZjsDzAXE1xF2tPXnzh7d5LfwYXJOdz0FgIDuVm09Ubw38gXmzTVte
MWG6eyjxZXnMMMjXhM4xyEhpmTguT4qaWBG2/TacG8ITnG8ULJzQARMqVtLf1HsvNvdeJQljt20L
dV8qZQCG56nwTw7qmJQ4k1YuRS0EuwRCA8BezbfLJu+sqRcfji4sDa+aJ15w/SwapxbvC/LZ45Fd
/CknKyg78J1FMdiIc/WFCFmj2ukCCUQutFG45cFWBuDtCqapU8vwGz/1MNmgX8zrsSQir0RlR8cq
WqFRLCH3z+Z1D/zMQe74+/LgfwVLPgGBHFjHZ0Pa4p3ubeGi/PHYqetmFi328OF/btv0w13oNYn5
/FnrTdBz+0UEds1LfPp39YxXt2WQKcaB8At/iYw14CGQFN9YhbHSrXN7JuhtD5j60i35kxqqOmSf
gpJEPMH4/WkLBLiTToEuonH6vapGLo6GseJT/Cf7V6YMnkuPTO/lGS9BmPtyZVyROMaghERkkbSa
PXP0JVQ05wWoYoda7dKPDVk6Mlv8omN6Nnc6FrPxPpHiHHgJGv+fGWfXMqE0jS6yw7/p8YT7naCV
IIaULTuEfDc++aJ+CQAxvqMFudFZiKBlcMjKKiAC5bnpf4ssZhYMShimqeuHul6BWGmfrIxNPTIG
gMQ4nPIPlgpZD2TA/ObETBrri1bI0Ru4Prv3EirjT5bZquWef46rZTgOSnplB8qMp3rHJnoSAS+o
v0gFze8VPvjfPMxyKEvW9kcd4dP85JyvdITf/BubQFH+sfxzaYMH6r8v/QlJ54QoKYrbyQeqhoLp
Lr22gperucUO+2paxvZ/k1mqK+O4Rh9C7wmQGmTqfXXLruS85q3bBKe2a5jmpPy4r9NgIEtpq+Ae
og4JPmdoQzfId6ZFlGpc8Yj8IOgIb+tKnjt+F27Pmq71/8ynakAi2Z9D15cKddqFYawQiBQja5ff
bQ8LtH9zSDs0awjGP6Q/O2cQF1fdcYqroiyRIRU2SVRy9DfsnHGtNzd7tOONPb1SquUIvo4OEobH
ZZ/LS/w1/nRoFOXI3AW9YHWWKTCbizLwUUoi6N19coHfvrQ1cLtlKhndQ9XU04FiKbUbncwxuj9K
auP3SNg9O8wLF87E6SKY0HxXJYYeEA0slcLGToQoGh/m393T457np9Q8gQgBnm/iIp6AlIAPKN9o
RZ4EpKviC9CT+qYOeBrOfckwZBnlZEyckzd/feIAnYY6yNc5M1cqheYp4Mjl27LpKHC+BYfYQ08f
8DPffQEmCYFreo8TSk1pOJ80FISH4ERH2MXmRmXr0AmDB1FfP7DmOj7oGrI+kAxN/mD4x68xFouC
eJpSf9Vv1LrOj/ylZdWKGIBatXfhkzUCsVDku3Xm9wC9T5bcwkrqLcS35yqtFK9fvU4HomWOHwn2
Az2I/GGC3s3wtZP9Jx5/+KyjubzgI4JdwSLSJIGJr6jInJ+OnH2MrdugkE9bRc2wJOKQvVsadqLe
BfqEVub2FADy6jBLqQMmXEL3hBmJDLJkdc6qwZJ5BSur4ysAVk0p/4gQSbwI793xqM04fRwmXf+T
6QEWAPvfjIGcOtG286XkrQwukIhFW7v8X6McuouJQ/0BkP2RT5mbNay2W3ifs4Ah1nk/9go3f3mA
LvDv4i6MpQNbAksFY0qsEgTp4HIZoPnEvoqk/ZhgaBiFKGioUnIWtWm4y4aCZUWqKfp4UWd5cL81
4J6tS8HIY8D61Lkud4BNXrZeVdkU6Sf3VfPvRuNvSWS+uoblyK28xeyIJZNCIrKfBMP3ksamMLp6
lNfR9SezZan9NP3SL00fBWtfL/wbuve02K69DE4tMMb4BmNLkXBCfx4qGGLVtkS/EEGB8RVf1tWX
b/zfPrbY0QEMaBdvEHbbSYDZgOr86ii/SurNtnSAWiLB28h0paF+xhG4G944ANEMT4o3p70rD5u4
GDe4ugDsY4U59r0S4kXgZpThQtI3kUaczs1H7mfZQdMc7QMBo/pt9+ZSfuhFvyNgkEN1FD9KX5Vq
pp3VsY9VV5F78RaxZZXi0/RW18fnnTg3ah/XxUCouid7DnE8evbE/IUzK1gVVmaDsSTY+jdQgQKR
Hyj/Zypg1Rp738jCQq+p/hhYbZKPePWnGXzDRPhdXY2xPz4J28TqzWoi08TitZGRZFuW0+JUR9OW
umbh02KkviiuKj0WWIEtKKjnRe7HtxNSTbfInBdyDfundgLNvX9FUNcIge8ZMD2VEXtUlmQ2BE/F
ApoeFosBRKOCjgTQKSRXRvblclm4nP+paJ42pkrVEi9vDzwEZ1Yx3gY0fBufyBEd6MsH9XpFMMBB
QqS63F5mwPEf9gVbLqhSaLtiBX5O8mlb+B1ohhLLBnujitu3qPCN7pMBWfwYulDFD4RmZipqCAWk
xQcxKF6gbJSegmryIXWXbwx5xWl8S+b3+bCaIpGdyN0d6L8eXQQPvLwrCWd/NKt/IpWd9PtDJRv5
YSwinAEMa0cimRGiO6Z72udT73eokFaSjtRFp8EOByxE+L7oLkmBY+7+DFJMrhqwt+2DzjEAuY+v
8/IbaISSE+f43VnCAIw2VxORMo+UBG9+pizvOWTHsroGu2PW0zGMdTD9t7vV4NKywQbzs/Sf42da
KVfoCwEuJGB1RwXJxXyFoAfBlpOs1Zrk6oj/A3MTM2EJvNCKkUMJjzBiYj+Ek5PuPD/gseM6dCQ3
OW3gN3KZNcCVvVkNBStE6QeVN7UuNwnWzHN/BJw/ztQ3WC0YKlmwTzLRc1zOTsR+0o3ESo5ee/Il
jikQPX24DAOhP/Q6OGBoSY1QzbAY0cACp2n5qooTx8153yiJA0jEwSoOxhw8qpspOUysoblajXZs
/NMAXYAtuQboKeD6J2Oyo46lOic+mGQMStEj2sO5CxnRv23R/o1BHavk1O+bbYeNcZTx92sVSj0M
EQejVli1oPOa1/eULRPXSQx6cakdpzqMfMa6Va0L8zlogLtr2xn47sxQywCQ+eVsEVDg6z9jUOJl
NYCKHAlZfFG8zbofVaI7q644zWFIObTbgNLzzMuWiPJv+uZ+xi9D7BXXJP+9rT68BWhShNomcURM
KlOGahiXy787wm7E1Jg7EZUc51m+8LzYZWN1BgDr/BZVcg2q/b4SJ6vuj2zKl9XEUlvqeTYaDfpm
gZs9BKgXjeo7c0Nv1SZK2Z6p5fjpjVCk52iU+HcZvNkuSz0XmaX7s0dZZErM56/FGEBQQBwbnPl3
Xyba3sbZJRo2LE7Yazpfs4jduhy54vkBt0NScBy3FX0jLt86ln+yDoYhCyd7doonly2l9cVIFXOz
68Infu8kSRsJLRApNAE8LnQbBfA3x5DcR1SOS1YIOpgnJP/v9uc32mWh9CFS1tjX9qKvBmHh14le
6D2z0A3Hv5U/1/mNBwNJjt5dmuf3WukmXLREbOVDYb3jU1kgDvgm4qCtdw+L7TvjyXTvVf9c0Np5
MawE7QcIBvCk3H4HpvnS9+xTV6Il2MIAfdYtXphDNr1LiGWG8tEuigoVQRnuyBqPeAp/0V8ZjDOQ
SdU/pHiQn3dxwAp2khVkl7aqEu8M9OHRiN0JajCBPjX8qk+B8oYGvGDl/Su6wBVoNbdekQogxJMP
RYi79UHWVnScXf2VTnbxeqZswpNege7Dqa1HjnjL394krrdV15F2dnntDob5SqpkVgMKPEBOkDly
kqR5WRZfq6dqn78Ibgk9jROr/CjcrhFKbE051hHTs3E8xxZtYkdgEp+Ys+xeGepipvagfbLTXisD
Y2Z+L0UpKFmfJ9kQdeX/62kFvKja2NszZBY8F3FCU1xjF6jBe8DaZvcPkbc92n/w8fBgrq2VFRA7
Wn7VH32x5J3CCyzdiXW0fqR8AHHKJCo7Z3BzoHyPOBMckU6NxLScPBRCKLiU3Y/rhx4R5VT/3e5t
KUQSna6YOpISyNyT7ET8E4NHvFsD0AKmd5z9+PkGk34bBThVeh2HH3ZlXK5esJ3G6zRgA4jcDGGD
FzQhzOb+QZ7UtZaxpbAJb8GNSiJUTZ5ULu5k1ZFVHL97vi37xV/PZ5gxM3xekjOzg7tKYaq2BnWH
wLkAjJiTZ3SIpGO9Zrotm9br8NQvTX0em8wNUL+VfH0InXbLJuWLm8PUSfqLEqA8dyXEcZmy+4K+
TjKwYlSjbzeVz5Eo8DJdmgPoIz44MnJ4Q3K2C5Ox/T1+1P586K03WYY/54+Zn5TPNy6cXzjeH2nr
zU5YgvBuNY32j2Sg4j7pB7c4tfDpgJyOdJVDVBv99vNEFCbgjMf23vgqxf7HNXtVbdJdK52ls8gk
fOHhbIMb+Qskoa094JMQK/5llHtItBTXI5npq+lY8J2x54QeY2U+J0/6sPmac/R1ONxLN+Vj8d50
BuR5qzeoQ0cUCE631Mbq2r4YMHbHm4tbie8HO4x0/2hPsVlAiNRHR3ZCwIAMzugDNiOVuoD+BjMn
7aT8AL2IPrUwBKQUY13oL3hpa1dmi0Ex8kQIaPD9lEbVyJ95wb/WBpVKMH5h2+TTn7E5/pHnIBAG
I+GSoYrpjXzvb2co1tmgH0kzyVqOjAwVFhzPEOIUkYInGFJrCSFnbCsZ1i4YyCMP1gnji8dv/CZU
g1khlChGG9Ap6VTJJGRU31qAYbCpsaws3WUrqBJJTfvlL9MMtWNR+TSg+QzsKE5cOQDO4VUh8rf9
bK7ZtF/AQ9SeI7vZs4qB3Gb5YDqjyVVY1f+w7wVu2SpECaE/uXdf9EseeksfD5xmV1397aiXPn91
0Hm0blbjv6Yw96chWSH+qS/L1ag352CvM9ysty0CWfcY6e6oAA8Q0VXrrpvU+TE6lyo1+2gGvTF6
Ui97DNZM7txGx8xia+AhbZXRnLkqf0yVXqWEbNwDo9Upc8Y3gRg94OI+xa8MTb5nYOyFHQ7oWPVD
vWDsMVAM7NI6RaW3r4/+S7JygX9D/LCI/cjgLZ8qGAeUwflnLAqDnvu2dHtCr4834QVwPVnTiJzp
+1MAC0bLNChT9GWomlscHOX3r8nJcnwn8O0Bgkt4vRFAWBH8B4cDWu66HHwXEaZKpt3nzhZbCXLW
BV1CfL6p8EFSOMXp+FUVmPglORaXilQXLqWGxPZZLVZBw/Zc41x+gXXbOh67GDYtPtLk/V6l7awC
c6OBosMoKKTm4YdECO4hIFUhmUECfpSMvr8foIf1kxxvP5NBXfE9MnYIEOfsaIYkKrEHQYxdV4FL
1cFiZa7glFVTOw/66Zn6PDuo7FEQJokaHiH4GGia73LxmTrm9v7RfoYMGnVHxD2jDcMRkl1lZ/g/
ZNoMOXBSK6qoMXEPyOOBDrIOUlC61IZcKmRxbx9RjVA0VkCGy9vY6mS/Euf92fPT6fTQ41wfL08K
L3UZxc4X+vf5nEzFSz8oN4XJERng55WaXma3OeLrAddroVWOCahqDn2gcT46684cWZjvURXnfOyo
oKgE/uTAFnSebUhohY19xUeZiJzuGxdEeMr6ktXAcUanUSCuQjwYc7vpaXlOEd9oQHlfpQ/G5ASr
ZNNDjnC7DS8Bz/JB8uGpoKSbKYpDe7H8AK1E2hogLN8wIpsS/71MvRz4ow8YCcRa2HWBxvlqeDvT
k0GuATl4JV2UvpYWzbihbDMn5xbu1XaaDvw73c2OYdeqFK1IJJTND0ECtk2zV5kXEo6VX6DrlvU+
EX29dSZpkzXEWkkSA6fBJKU1sAG+9AZG5KwBXMGfND4GgtoN50ZHgkOtjxh+NXKoVvcgFntW/TNx
wytLPRAdDUWt5mi2IJZfe1cYiNPS+T6+cqjS5Gc+kLTLCS5bejK6JZX936UhHNQWf9NZIqeDfzPC
doKi4sdIrAlcvTs8xGoAU1vbVidrjujGmYjv3aZMnLkmG6u5OkohYunRg0Jntvj+E7KiRvQyVE9R
pLiIFjC/r2tVmliSP3602vBBRtBRp+eRaAH92L1+9CTrQ5st/eUbkpMLp4uzJWLpBEjdVBeRh19E
2+/W+PVgWO00WfJoKhCjGI2PXX0td+B0XAnT5q+OdgLVoLz4mKE9RHNtV0G6sc+jXGEsGtevCFgK
g+qoKmeKdLDpGbjzpMyiVryCGdBAW1GctwtpwcY1gW/ZBcSUWP2JbO66drJUlKIpY8T2G73QFn0J
JtD6PF9l59vmDUjXQ0+XEOmsYuOYRTp3A31Exc+KD0shMN/RKNCHeJKwG+0f7/NM0Ulksb5d+NCP
HhGL/PYqGCPBwjn3sNW0maiElSJ3hDfGzY1Ab1yqcKRAgrEkISooByNmRQIraYmN22VC/MzdWDoC
EVqBSSGSm7ygC2ePRIPCgRR6PDaQt/JMs3t+7NfQS8Ro16m/VJJQpfMvr2vHrPhiU5IVQW1G5nfl
o3O4Bf4/xbmKScWVZoUsN4fcqd06+XMFgeGiwed/IpMWSK3E60fzj2ZIyazqf+LDLJ/qmHiXb7L9
ajGBcu97yss4WM3rSfNzeVoOaEDHrs3NCErlcs3T4a1nX5OUH1Ma6ymk7Eu70Y2mM42YOwsGqoep
k0tKiKXgLchzOtQ6E4bE3fQXooUYdGFeNAR/xUhhosQtRv0vDp5WF+rE6FWl/F2wi1Et6uQG2naN
nIt8RIgd5ZGc9x4EV0DBRjUElPjO5SlfPQmXQpAcYdg4+GdaOSJ8ECaO12zxRbB1P270PYRol3Ro
Z34i+ZCp6CzCgvjRivlhVk+VpIRwRdL8UJPCWd43KUltBvIoxbb2u9rBsk/aBK8JoRaoma5ptSh/
geEaivEpQElwBmpo8czxLd1IT7FdssIhggXHv54slHLsObrwu6BwFfNrkv3fZJ58Q/MEJxFZ61th
3DWTOklZhhFZuncRNJPUOBFhmcUgCY2yOK9IyZfbZJZ5mFkhqSj9svO3dxE4+txLE6+sg7gfJd+E
7cjQHzbg8YsjneYLYtnse5k7yTG1ajpSF/DEVZYmRhh/2xmla5hFehZKxqqRexvtIpQ85oN+ZfxV
RZgH2+zi4msPVb4slZ/ZdDwh4WuBa+UP4dOritWO9k5+kNUdq7fkyRGIbWq48jAHJCa6sI1eDWRl
MrIoIPzaPsqiAmfgIPgUERMBVYibdu9MSCWY9PeqBFxztG87ozxlWaKGrT+sHCijzOKuVbgklWt7
evFzZ2lh9WljVJsCB4U7FUmuLfardr/0X+J2anuELerF5nv6ryuVgaih10nU+geIQQB9L6qjEK0R
pS2NQDUvAtPzD0JqLOZXsJBpbNo9eSPJAPCx8eFmN2rveBxrR7oc+Jc4enAbP/nQHyMn43zAWUC+
I23/ErRFm656+SZqlUzXkmm7TqyanMAQEyk1Sor7F/lNfnhogaFg+yMA/G/V1rzMHIjzO2esWGf7
FdUmpPy5G2/FDCTRZZorFq4F40kgQ0QSjggM9giG51u3yv6DuLjSJ7JGF5SQVN5gj0zfCbvxheDh
J4KYQsFoq/rOdY62TWw6oNkB1woWDZgafS+CwYDtxIHI8tKVJPQ42eRamMZduC34IQ0kuD2pLDIL
cjtnh5Iatpc5rZQUgZ6yAQ5THFXx0IFxj23vJLQIGwmk7N0dVJ2cz7sZFisXVcl+AcGbxEhQJks1
yxuyEc3HGImD18H8zEua3JSMGZPDdVHCWiQ2WpBN00tM1U1FwaQB4yV3iRg7EUm3D8nANgmsXB2/
sjrlHbz33WzUhUFcyhgzFNtRDOTi7mhONXqXuX2AJQgQm+BTZMmcMbOeKIPbfqAf18WRAROfva/S
CFmyhWGQPsd7PtrVdD4h71N2gYRwaMMhiHna2wHGxSD7BohPORdeM0mPAZcAvB2tmKLR90aZorZR
6B5I6gTot87ENR3AbZ+GomZBoqWPZmkXwN68H+QwFSsS/sYqE0nnO+ppALcISk+xD+5+xSR7d68W
o3L+pBSDY27UFz+kbBCXUcL88mSdtyTQruqjNevw44D0ONjyi8FwES5eXS7krl7Ima5oZWujUpre
0CMsEn7wD+vCXj3/AhWISiiLKmfyHvBWBVBDkI3ao/rKv9Ib6u/SCC07bDAGFMh92S0+kJ+2R0I8
bc3Ow335rhgErfUYM6EG/uRFr2QEu3b2jNgR8ExW8/antXJ5QK0nAR4okJdfjjUcyxTuOc8niWrW
ohIk2/by8DvJAxr49wUaZLldYtxvqzUorl8Ghul7AgO3H2W6d3TdPyVZd+WRLrkQpomxJAtAMQoR
JsXgo+0CvscbJzi35pV9NGZL6NqBH257dpn9/TWdgQE/zeudX92RzuENqmy7KkoSkozu6qF38eLW
tjsmmU2If0M2OkjhIghC2qM3Z13ReqGKIlrpAzmO7GgWF+wQj9tNsPUGFRavZPNZxdPVmTu7DZVt
UTyrACiGW7rTBSP6o6SilUZQmfAykLctFJrbUoAMpRLnLojyWSBwHWUhvAxQ1jWIu6l2Sr7qMLsy
8pyGk0Z2K3zkft8gVdR4lxGXzVWrYLJ3/8eOer4pGv7tVarVyzrZuMghxrV8Z3uq0lhOCWO7Diuc
dwjGdjPlVwfBOAOIrp4ErVnf19VfLdUT95oemshp+ZBpqI8TpYu30G/yJVa79svRBFAm5b4ftZyB
gM7bcPgELVL3iZ7IUG4KRrCUWXHzZYFi2pTRGSY0fUIoJC8SYJUOqZS/pLpLpHQC9Y0586MtpDSt
rZSi4HjV1m4SgCEK1C+rdW+YAF+sHEZzqUYUG+g6fZyxzG16/XpXiRAk9RVDYpIj38iyONTn60KR
8DSh2ymrW9FWO4gAwrTKc/wnl7fJ4yksfoLZAPwdYQ6RAX6IrBT09Cra8aDTXxH1zRqVU9Npj7oA
zFz/SIff5IdPz7OPuFPUaIGGM9Bt3ZlVpNJQi/Hv5pvk7gXTNdo3WMyA/IHeviXwxtx4ra8uYHCQ
+h6grr7S8kUixQy1AwIjq4sF+Zfzr3oEA9k5qm3JiUgJwGHVAmBN/VDy7i6EZqX3Fj69o1eHjh2h
c5PLT0PuoOlXF1KzCG/16emsGZU5bNBGHa7VkOFL/mrOGCcPcSh5VgsYaXz+fJFWC4XkYBrsqTwc
e3Bj3W11PPglaKJpeTbp60YHP77LCVzHYjh3zFs9tlzBBZnysn2n5zBO1qq0QrdcNqU1aUCFmAP8
9kEGrCbw0AbkVSIhS78p1HVzSSGZe8x9ziVx1ds3kAesQhZVDJVwuv6hQ7ONufEIZDc7zS+0LEhr
GCUgL9shAae54X7xcussbeprqxBtIhqC2v2RhglPqJmscvUSDYCKDTfy94OkJAoaVEtHuhdVoaU3
YnT3TphYnj1EjZP7yuE9IqB7ulafMgk8DtCoXftJx4q2lo4P0p+kH0w053rBRc2/BoMGobkUhx4D
f4XUPwhQsyAWDesQNNMk8kyccFdbTvnRIhFmlKI6XWgQqjKlOxbj2kVSYVKh3m2l145Sp+69A/iu
uI2dDk8/1oUWuTMMOo3NzGMPTuVX4qQHtPPJ1NMrMt3K/X/1F3rMHXYJZiBw3t2rqu6T2Y6EJFfV
QsxIGHLXlSTjp8WnD9hdkzvvA2x7NyXBAgfnUiR/+OWmk0H9Z71R2s/bWjZvdZ7XaxHSm8dFJlJe
K+U1XRftgNTIPJniiEka6PlHP+XKMVJ1ooLfJYbzvnclbS0mcb+5Oajf9LzBQXW+miB3DAzwaowB
oRT8/Woh10vKlzx/GYbjUmDvBqqHJt0zLDd3QItCwf4QIm4IdvzfyQS5XK+PF53Fazw0iUBY0KDE
EFbytE6yN/aUPnLmCFlxO85HK3S9r2keksWBNEVgPRrpZdoctCKzoRBgWn+Q1FU7fD1judRatnDe
i7OnoOe3sKYsrBbPgLaWwpCQLs+78tIMbLEB8gdibYZnd48ANi7DiLP64Jb2U+RPSXe15IPEx3X9
R1X4lZyvWMchGqMy1uNzstfBUIaTvgs8luBUPUWfNBYCZuSAF3lal6SGoi0uK/xHYHMs2sIRekCS
e334sUTN3ReiHWqYyHyvNl22/lvgP92gjphMGR3vOW1ht7b4+OXy4CEzSI9PnB7DsnkM7jYCrxxW
RBUoNw4SNJM3KOkSFcFAyylyiaKFCOTaghYB5Hcx6ViMieKPEa+V/0tWz0cT4Lgj6YyZcXVCwCu1
O9sHE234c3f7yD2wdjw6pV4uMNR1v87YdKK1tLaRRo0nRUFHjAVHooovlY0ytU0rYkrujJ+TbN4u
OgYt0Sxcuk0IJTqlC2r4RarLz6aNBvp7hXBLJ3VNZJB4dN5dHAlEFEX0sxJqa4gsBYjSOl86zwAJ
WMNfMLPsF4if6wDDd+GbncRFMdUGdBXEvdwjE5l+8V2+y4FyQH3hbJ80NSGGDHnYD9FzEY8XFsv7
pUB8+teuIq5dZ9oRgPgSIX73uaxpwo+zPfG6Lfh8fIulaq69bVP8Lxtv7xD/mFGwha+HulLvEZ1+
7BpoQNYVSvNZBcPa8T0Htazn2Mmqs8YA2Q0WW8xlC7wPSV/G0B8pe7Qjz3SMpB6YaJi3DqDCED7F
ol5GJrGUehcA83tObnGNlV227r93QnhrngFrDg+yEmEWgn5yUtT+2Qb2/6wIf2RJbbqEIse6AFWm
fmUasKbTmYSnuwuFLHFxh4IGIpQ7NI78ZRpPRws8nubZbkhTTI7mcjgbPiTAGkIQtE0BgwjKrqPf
bzF4e0E2MfsO4U11edYpZawPWJcA46Gdg1b0H66egxKDfGhV1Z6zGq4qm462KDhoLCSoqmqh5/c6
8cN9wCQnlkbOUb7TULI1jtbce8kfcgjkOeiEeMSKb7VZJRj/+ebSAqEeN5bWIsAD8QusdiRz1FEh
7+NlZEVvUJBhdaebx3QZo1kVA8RlTQe8fjSLFypaTc1cW8pHJfbspeCpvcrQuPGrK07mqOXVFCHe
EUiLml33T5nOyp5ogi31QwtzQkZD10vMvG10sBY6Aihf6MZtmYAuiOGrj5VgjFFR2mgu4ZylVoG5
IVL5h1rCGm/elEf3YvQynS14HCutQa7P88fmqqYolMgg8Na4Hb+VNUqtA86QEtapYr/qxIOHO/NH
ES30tkv6U0Oj0ruQ/o6+16OXRZm3Ie0IH1cZrB/3VYtdCvOrny3qBLbOmfzYf5EVVbAFnP3dbdgf
Ri7NvLpWOimmuH2gTr7e1NAUtFBagoHWccxRugCy6ZHiqyNgiFoZGrhYYGh4NTjErTBQn+w2vSRm
1G2xFb/ELdhpQCcxY066ufGUQ+Uxpym6AzevJqOKUPdl6fbX6pQZ4dAN1q1RrBniEzfaxtCUU8EY
1Poz6T4aYv6ExV//PMmHhGKo7VVmwRieUxJEoBEa0KH+W5PJnfo3hRLjmY7Ok6ffRcP1yw4C7AGF
rJB85yAGVtV3mCD8wpbyjgz8eNADmsPelUObDYOnYFiPB3Hnp1IOWH2U2GUwJp3czxu/HLZEBj/a
94po+5z9HqWOVlw56Cj4M6MI2itd/jIciTF5KcEPN23qZU3p4G2FAR8QJJFzBnUYTMq+PGMauQln
3fOEnV3hMlbDDYcqx6JF10KZtjqQODz+gwt5eGHM4vFjRjrxp3FNGpmzZ7lUofeldTvpYkFv6jRv
m7bEbSRX7ae34vKdBTiAp7tjNOdkWt0ThBUSAcc6IPeCu1HjzD08pobV8T04Fx4N7dK9dB9n14FU
J77KppmoL4pYLRk4QjllCLoz9VzvjvnA1cPA9Y88ZEFfUqZhvc/oU+RbenkvTFExnxd8GBYewJC7
+Y1kFl6q7SPkecHmhsCP8uDnL+iHLhqmUtiaQ2vRGRA0H08A6LdUYUdSs37RUoih1mG4kYOmyOdR
jWRvUc2KpVPaBDKjmtfeVCMr1FGX3Ik3EZPV7gaJOmV5/hWD7XSxI+VH+nz0NYa64pd5u/kXpVdD
VIBjwn/YYjA3mOfXUOtzTcwBbpbl8xK3pM2X52oB3xNdeSamRjxnyUMDSEoUSnUVxzTp4P4F4whk
1Ch7/sM1M0JFdI6oBu1IKFyydli/5VDWFbP4Bzdh78wKXju6hMoCzhmS/NU3Yhe0eoqdGCCzbANh
Ho7UkDZksLxgA74d+UD3pTdu+2VILeY8b0XQk66qbcrBwlqEe5frnJBrY67thZ93Q+Z2PPVe4v9E
iYe4bFIMXIITZGNUexx/wl+i/pGDEe55TiL8F5KtHvnhnR8WXs5IhybrmejtrCt8n+fl3a339OkV
aPqU8xhbuarVCGZXjYCoRKTyn1MiV6paU3N0Gs7Ze3TlSzxNPgfXqRQ8Wzy+DEaFUFLq1oM/uaga
msbCRf3TQJpd5hKGUMut25vwbqaEdyJVkFMmoFUmERKwWnGTc7y7nXFmpx8MdwE9GaoX/OhZcLPK
6CKJIH1TcTWkQyvUBHQLcMKjr2qQuJhBvp8DGLDs01tkwapC2zCVpIyxuy6FyGKC2OPA0p5KLY6R
GWDZpzpNwuJ8hyM84ZmO7KvcKp9Sb+LBQwyVrkxEqi5JsD1otLPDx7lmgTvAlJCPqArTQFoLAD63
tLU2amA8c/LwlKDa2JC7rpihANr609mY5020HbFuqMfQ0CfhronXqv8KyqA+X8MT/xnodNAyI/uf
BMUY1P52QMAFWJzZuzk1QAuJ3VabmQ4cgy7hZSKXZ88NvoyFEYOeLqYgP1H+YulBm8KLpaAizAPi
u5cKAX9vxuImVsF+5pjMMOVszUmEg56NBKcrkXg8Z2gjoXWXA8U1eaiBRkiYok7XNpAb1Vrgd68w
vtU70fpKSevxIgnYWuQhDblZfBVM28wXYlUy8xeBZizmUQ74o1bsx9ou9sXjFWtjFOstAVotqCcP
sMMYi3o/50jCqYCrC2oQv+K+v5G2ioFuBNcNj2Cy8Gpix/OsO7+swjvJyVTWoWqZMhpkmKj0L1E8
7mpC+Bo2erdzwixdh0oNV+oAmhONvVANKgp8j68ut42xVuS+6N/8OsJ8Q5eJk48JXsZwvm6JUeuT
N5jQMCUnHiGj6G3ElOBHJZyBzlGhps4CNZHGc3Kg6H0rupl4zcvNcyzj/KfY9VbQusvBCskY6f4l
SwZ4wBG2bOyxeY+rMqANZ1l25Efy2Z/uAPumbJWPeXKzBxe9u6ZVRXP98imLnRw6z2Kgew2FMafH
URT9D7Z9kGoU81B5eUhD3oxPTJ9kNtySf7hwIf3gJINsW7ZNQPKKpIMFveyYjhL7TH6cqRJmVyJ3
ZsO4mkgx9keXfpm0hAMD4MOjzH777R1oRnxRh/UNEWUdVvkGsU7YrbYbVh+WVYJ1pm/MJ1YIajZk
/0xsrXw7O8V1b6V8saxbB/MDrjX4zFJUl/I2oqpqd7R2hHU/Ncg8F0dE/NfjW+6kTzEJUbE1uBdS
xpaT/NHjrmTHLbIxDjyorrE6PMxBEJNzopGxdBlDV/h3K8dGTfC3WsJsSbRclzz50aD3ssnKISan
/Nnso2vTqSpSq3QBvu+pTgBxhmXHo5F5fuzespmi9UzdeBOr3LxyeqeOd9uiqBEoBk3VkFOHnOyB
2AAr8C7q/5NMUv5xEuULQr7G0a4X0THSjecepGmOTkohXG0fvntA2WvsOEWad58c9uAyXwTuFFfF
/qjiSvpWA+dDxjJV5xEKxk+JLVjf/MMfqJnXael2qVNbifiMsSoh778eJhgCARV/3MNHR5sXjqLG
HX2D//N8WwYPJI+GkPgQaHX9bet0EqFdKfP5AHKHLhzm+8dkxjHxfD37Vkej33Cpww7Kbrnaf8lq
ODrtH3H5+jIvAxpnnGJH4dbO4P2Xuzs9NMbpJg5MPm4YN5CNyUFLckdHlnF1x60ZCP2Xlq+4KjfB
VpFYe2UT3Uiqv8aq3AUMM6U3UQ3qlUkMBCvRCwjMyG7c9wgEe20LYyJmLaN4PxFrRouf4tGatLyq
tu/cEvJ72KM/fH51qYbjV4vvpwnsGECXu2oChR66pW7yzrsSyMmYcadozV7UK1y4DyrXX00L9roc
ukR00lKeqy1ewAOVdthsENYU9DA203I3d1xZE1jS9BoyzlQqGtyAkrRFdYhJlakSuDiQ/YqXeGM2
JAGvKHZ7BV5EOVd/y79MItf1pr3WKuN92F2M5fU9fePIJCoGzgiQjHEbm4amelo2JMPEiXOWFZhU
qYM9wWNidekcHZ5fBGMDnq6XntwQSdI7m0j3s03aPTMbKZnMJmWLAop2JzE0HRQic/l3+xsUFrVj
SI1D8MQlXes9Lr4RWUP49fhNRYlHVhxuOSuim/nbptnlqgjksA5VVbILKX9Yp9/8wbl/zZ8X+OHi
HU4ZgTRu76hg2yxyjKvbmmG/MXH13hlV3BfRRL5TAmyxrlo25tjPkXHYKJ9RUVCcWkEKhxH1An8k
e2mBRdY+Dz56h0SFlbjH5GbCGtB5Tb61GRSRjY3xovQj9nO7CmBq3rRLRki6lx9SEb2tHLeerBo1
ByjuXbpuE5P9cTF+RUOiflmC0ETkN696SBWI1rlnFkBROseAux42E2u0PCrfP+pg+GRfhXFMehJS
Yhr5HfaPGUAD6BcvN+v/Y8AEVjQbZI/wYTxXX3eJFdkMG2E8odbFWQqbRlMzv4zMaNFssFknZTIE
hS0WjJKuv9FbhxlFihQ2w1pWzw5iUZDO2w6WghqcxMrW0uUt2jm6zsTenAlia05U3GF6XiP9evGa
+/wGm40JN3ZTUMBZBPFgF3i4s5N/EKWXBFP1fL/qcQy+H0ufZB7kicRT/6rpHsGhJhmR1ZG2vGVq
u0L2FF6Mq4cUeDFItp9eTwl4+BaZKN4kl7FKZLvviq1OApJncOJy+WHtnyc80tOmJiguIbnDo4pt
9aetkobJ6JUPBrAqOATaiCHPwLzGSRnXbf8sUZ5mpqfTSrjFf8YUhwvw3ipMKoC32EuymWrJpPFV
fauSkIn7pf2DN4xx2AHgDEp/tF1irhCrC16aOEWUEcY9wtBv8UJOt1vCi2pSV2cPXmCZETC5P1kK
0dXdQ09c/I6ivB2i/At3E2htrL0NRYeHnRcTTXd8TKhXW7mNgX17UFkmyFCbygYH6UACGfngeCQE
E4OfBbv/7gBLayJHD6HoVUBkzfAwIYXDR5nr97Sn14cE7+GAVt5V9dThIDKwa0QUJc2zt+qRLov8
btQ1xIIqpMJNo+yIXYbnZpv91IDY3oWF019Z0WkPmQ5Tmt6LE5lHVxav879kXPBsymN6NktF9kl7
zEV4lDgAP71QSwrBQMWTvyHpXjHZ7AblYxQ9ypSg2vom+ldxwU2H5OQA2dMW1AEwx3EPHMr7KTzs
qVK53XOcLpX0FIq8RGDqBY7TH2rQ6dOWasUNv/NRsM+l9nvzRHhrwRC9AxlO8SlKa+oIx6pL9mjm
gPGXTf/3msnk2F7tJ0RyJR6gIXSLk3XCs1zt0BP+9JKRlNA3WpmoXxi5aZznBphBRLc2GnIyb+Ap
GcRNBOAbx8bYXqIxWsljOBDAZxDoDvp8I7cz3YUJOQiu5EVnmlNJnT1mu5thFv8oAx/SjVFaxwi/
2KJfCrzN4l7bFL+bkyKTNmV2cq6QHqsq60WMOigndqQyC0GY+13MpcBJ+13Z8lywok0lRpdQMuqD
rCgxv0Q8BVfaPtNLMWvGhmHmpFyofY2PSa7Qer1KQfqF1IvLy4AK2CjXOhH+nClU9UPUizhpAjty
/O3A6LqJ1UFhO66+lI3HECz6Xzgsa7K6Ov6MtkQUPld/v9CXMb044bjpRzomr+iQX5RYedMISudU
Y5h+X8HHBxGaOSunHiVsc5yik5ohBzV20jyDEQfFB5xxTUnzT+wQGGkpz/MtvqnXcJax4XY9oxtH
qlPCr6Jcq8FVJndXngqJScH1u4nwWsSOENK4nBdOczXU5+JfbBejYBvoFdAt30XiWDXrjzB5ibBv
dpBFYD2zhf2T50sOISuGQnbqaKiP5oIJM2iRL4s47V8iNxmotzpcBo+dLG+mAB28EXS9mkC+Sf5N
1VqU6+1uX0RLl9nhAN6syJnEa46H7nGsR58FkIvQMPHHuJGGuTN99E/xZqMZpVB//A5VWoMgk9kn
O/Tn7q1MfoqEIwljFCsfiykZslGE2ngqyKtq2jzMadyMCls/jdi+IY/D52PWAqKRM3+/Ju0nT9TM
V1kwV8DafRQMCrmbD77AWJYmNphawo5snMhwP2uBE0vbkC/qNgJn0GCA8A/gDHGl19LZk3scvnCe
ilMLOxWGF5yXNjhrRpmdRXbnanpM8rMyGGgP6h0cmCyb139M+DHgkwaqqYc691xMG2TyrbJSwDzU
hQGR95hieQM0eFWz3TQ/fqgmIKpYAQhHG0dCZPLgE2k+q9y1+sfG9qP/TIazOlWjFh2eiTKd9pmO
eZNFqugsPygrEd5SzeeQWNwAEloHS8Ey00DHvq2zc4cHgY7I7cWf/L6+b+XLiTHBPoQDNFHlpNrD
vlJawVxDNHq0ycjxaAu48an9PhG7x89uapo9T9WJfErcoZtLZm32cWoZrsDGsPdbeUsVwNXaTdM+
ErMcCGClyo/0LZ4Xf3IoHHClejfWtjvtUwh2ti8MCCNxCgtyZeV2SO0cnOXvXKjkTcwHvteOsMWI
k+INx/vPqhWO2lBdXeJqvEostgKURl3kTQnXUz5XJrLW2cRQog0Iepzr03luueMoaS1EDZCDfyRM
YbVXZVEL51IE/jezMM8zjJntjnWCqG2YaEOa/3M5Gs/imMlwtcHqqwdO6cHmaV29wzD9ds3KUS4d
ivVOT4MGWKjElsRevacui/HAlqsQuxe9fLukvxQy+3AoKOGs8KLi5SdElEBrR8Vg0cxIiFIm2rSZ
is6xJrBLXkDSIlc3UqYwiRDeehNOACYnvEPJNBqkbJ2Tr0jQYDF7omjUjElqXpSi76YQz9dKN9jl
4gDNsUWYiBQ6KHjogmTyix/qPG1eQaiFxc2GyYyXPtKKgtiuBg1MMJlJM4UEuiWJ/QeqEJKdzpxp
B53kuPrIOLclCE3yyESkNqnFijvpwKPCvuU5kCdOT40J6ohQK249PS3s8epcuv7BQTT7daPYL++g
tRwYPNo/GPA3voKAjzBHornXH/lmfoO128ligVDTpayiUcHO7aOG4OwxRGY5yzIcYF5qfz+0rzdx
PJ790ntait6ARL6ixor9M5mUdcNCXm1WJt85z+62/cTkePk4jtQmibbfiUT0+Vkq81W5d4xfa7QN
fyt/8okrYNO1CN7q9Qkuhw4XClpRiqC+ute2SRmYwiwO7UB9/L6bKSfviWvrYxjtPmz5ZvY94Bdx
ChfxCmy9o2ltWlsDCKqt2SJTUZaoLZPvKMcFotWroxX0wx00qew2XsgXPDwp3FWHveFv4MdwwJoa
W4DLqiLu+mqgErmpCeU5Mc/jhzh8UtPhi1mD8npQugVqkN884CtItUS0ftdaQfda6ddvuNiHknXI
4cue+oyJ6rmozKhBM+orx1BFgdTbI5or93wBDNYNuSN04Bn/W9cFNbLPAa0mY7aLrjh3exuAiNue
I4ZmkOiStXvhwGxxCuFo/BZ2O0pe3I/24y3XLCyXKj4DPKXGaNsUWjR+LarEf95CJ7oxWd0D1daA
QD5FZPhxbKLhEpwDZCPVYpormNy8Cvh1ZNuKp6hqdxJTbn/bQdlAOwIjka58JKO6tahQ7lPRTPTx
Ur0uWAlzExS1Jon0ZKq6G/ugwbES+dhJrKBikt68KA7RhJXEsCFBBOX8tkEQfQQ8g99DqQfIg096
/dE0M4VaX3wCFaPkaaJXqtdk+gYIG4We7SVKlFVV/qvQaIPSWw7QHwN5d2Y07wEcjnvBBFFRh8m0
Xbjv24mT9NJbl94zTarHntKABuvBf8dZYi1tv69xDkUpWd/OVCjGIXn/p+mp+oyLAvRfr3Ow+6bZ
KijIef37bzP5eMRzb4hapv9H4csszVidTITfa3u6vJYnMgkWBJ4wHxafa31LwMeduT//FiQF2r0I
LUA31ybwEZXaE1AbkgZ3SiLFSgftI6l58i5UsGLL/skVA1ClOcqHAQWapn6CUQehiH8XEU7vD0YI
TqRrFecCYBP2KGFzf9kpa89+YLMKeGnLaypSRxjTBvDmok3KYrh3XV/TNBcUIAlw2JZK2Nq1UfRy
b3HvRnWmIFVHEyCjhl5WtWliZo/tBLPB73yf7DoDBwDXmSv6wehncFDMXg6UC7z5B7UohizrouzX
wWgWdkpeYW4v7ZBeE6HyN8sEADx/hrzi7xF7PZZTxeU9wyuucJJpuPkqNuO8/IgiYFzwgVQrk/Qk
DOZ82iYTljOrFnrgrpn1sgiVRqsKoVgRQ8M3wtEs9KsPPEj/vf6zfg8yfAK/gnhjL84Jgyr6UG9q
yD1Tpcq42R7SG937SuV+x4EiWW36AlX+EW2jVGl516AXWpRIvzdVNuI3TYeoOE1g3T30BvRtYsTi
92PBnxoVT6PFhzR2ROJgDZb8dSV3cc6pV7ZGKN3sHBExTVSrM3TGZWGVaMOoeIxnoQYdqJ3WKksV
qPhPq9I9op5u9jQQT/KOXGhNosZmDIZ4gmMz22RBTg8aofZOG8qrMCVcI+Mia/pVadGsUv/zaOBg
/nHEbMaGFktpxrF4EXHiCEqlhfjSU/Ma+X6KBWyfUZDcCYk3qtHiXTSEuKmWH8QbpFcMT8arSrJb
Acv66xzWcHGDcYoKnMpwTGbpOXwfAe4kb1N1xbRBPSDl+61t3TNhSzc65mfUGvgQ+6tgXwgIMPYL
sYhyqiSNZIjWl42SPp8t0NFk8OEaOZVKEU2AOseVNJgcaeq+GhjEapUxAwuvRUROqwoAKAxb1KWx
dragTrK8EhaiDhK/ndYWf+zv7w6eE+mBsTgWWSZJgA+uQW9IX4mIaA9xEbAFv/8o1TwIcynZ+3GA
/bTUdTMBCDaphPNOWOBWlS+ELbflc+VtIRZzf6Wb4IRd0TLYgTrC1z79tNeH1UqLtF0Xa2YEsFlX
Z2LmWQoXcxD+8Zf0Su0qgbrJ3L/sIgUWJf7696mu7Ztqd/ibZc+CvRFeTV9zSGdJVgEGZ/ZeB27L
fHGQxGchsM6M7a3O7UKhq88zdv6tUaAYLhPzhO909UXY6clWlT4hL0giB1FxA/9kzp2eIb7aOQlR
vc334OVRJrw0HR9PsKjVjxWZkX+TKiYqoJNmOLL5t3fG4UChFpAM/gzLNM0g3gui7N3SCk5OJ6aG
4WW16r4r87ZMNTNSmtQB499agNnAE8eF/r/CfW/CxEWTWmmhSkxFRxvdKiXhOEpKrds7ed938dO9
/u3rpKKE+ogQO3zDUa9H8dMQx6HDe9s+8vr2QPf5uMcusccNJQrdF5nbWf3wb0ASThNglIXCpBxP
t/eA729+B6pdbWNEjcK5RZREzWSe7vXRxaFVlfxjndrmVjT94JCMRW+lNOZEKLRmzosQoRvFA8c2
cS9tLXG5XVveUz0hNcuZiFDC7Khq3QOlxnmzkhmu3Fs0rnWDrpS1klAO2H8KJ3tPnmMvrnbN3E5z
yFgtnpsNr70x43WfLuyFEGIF/iUvYdGHs09xnP3PMkT9qQ8onWiehySK4aPZOMkT/ZDiGlvX33v8
9V2fDDZHcPS3+Ceg/glfHdm91EygtVrGoqxDFXl//NcoBcY9l7IQY97/4nBitQ4xzLNL+Ol+NMXV
JXJp8P5FeeoY5iS/X4x4MQk0uGP2h5+TVSQ8EPagHK5XCn/8unEEuWSm7tuHwUtx3PadAkIE80a7
CG6KEbBlON6ahWLDynKscFKntB2Jf7NGPTHVjmPxkJzbptvfYBVZrEke8xBgTjmN4CgbYNEjqe38
EJGaHYb5K/Tj/WcVhCssL/yk1o3yBG/o/WpzgKk7fqj4SLzNiK3LvR4FJzMeiW7g5n2jLrkJzGS9
cwi+gQQW0uoQpFXgE0padW0hUc3LjZIlSyqwyApz6mBXP3hEP7h3uK6ApBtl6VGTl4moK83Jsn6J
ktRKXAnVJGmx9IwqG9ekd4T1hUnp+8gSqSbMg8pc3l/hcLDXaxkiT8/3e4SeGT3SUneebZ73hwaS
vQ2TKeY+XsPac0X/GyswVED4Jrfwpq+pG7y4QtJRf8pnMIeRmDvVH9qCp92hItCu0TiP6Pioo/QW
WFHgFa1Cm6KueEU+4fvO2iQImoMo4VM1SFEEjliaS+PeHvIMrFPhUO0D7KWS2UFVGtJ7pRG99THB
RYXcc1I3G98I2V8cZ9VpX2lJ1pu560ewhKFwrgqwJ7b7Bu9slCuIc6U2OBnljyVuCdoYNyxHSIS3
FM6um9bA9ZrHSxwtTd4as/5qxTKmt953WgFBMsRyISP2tCbRCbOsJpRIj+w7NYPSpMxPfbm86O6t
VYpORaCGQ8t9RTDnloM9pLejELNHRiJmC5juO75QapxC92KjC5BtenAs2iDeycB0XBQxicridqW8
1Ynt/tuPCDfVcaz0aEQ3+FX1/awufXnEY8ybmDo7vrAZYuUGU0t49OlJLlkJysTKoEAiGI3rMuBE
SYYOFBT6FnXX+Zs8OvCRim58gJZ9iHxY1D2qq8IGmFbKeYLecA64k+tagsIC/5Jv9d6PfvkLRyeh
ZeDJIKXs3gjbBad2I3DsPsWoHwaIEs1jo7vbGGrxiLuaPTfXWCI/07ZEXLWZC1mVIzkw+fJ09jGu
nvD3hPcnuUpbPf0Qdo416mOpX5TnS0o7uLOmyc/DAmsZVMNeVkFKxmmoGDPLpPNOEjFwc7E3N3n6
5PJ53oO7s4ZjTVva+uDg7elpFYBlz8/3IXilD4rhvWvzRUXhglsbH4T8lP0z07RC0Oi5Xe8nzwV3
S+NWpEZZlCy1xuuVHThZwf3sUD10azZIlwmXwqxuk5JvWLXR2xuhe5x6C9K3pyUSFHnaSWGhuLcr
QSmba/nJsrJlgQbd/eroFKux+ms7GaQ1M7Q1MGJkCISTXpR4Exx2xp00oP4QN5U792hjVagVBoIA
XoLBJ+Lf8GXV2YjWbZkYl5gX5VyFaXdeebGRbgZQt7/CHKp/QVOzllNzZyVVE4OMOiwb8dlrYR1o
awW5wkNxrqT8TGWT+Trx3JWKC+TyDc8DgLiICL8g3Q75tjJOtMt7nLLiwXti2HFialPV9B0WgIZ0
Eo6EqFSuTs7dqnziLZI92NVlm29zdQW9b8mie2EkHgreSJAwyViEhDi+4WLeLgPaRvtHAqJBtT0p
TccX/XWmME9iMDqKyidMGEIxQ/brl5pfO0QD97jC3SeZvFiXXDPAOjo0pCIpJ2tx9A/hqvlCAIia
o2Hr+WzStrp1y7nC7qcs9gtCtuo0XHfrzBvftDVWrtLRUS7eIadTSAVv10iPMctsD5oN59WzrUGc
mASdyEjEelWPO79+eUvhiy+606Oo0+7Olo1VpWInUs/omaLJogJH4p2tjAKxYBqib1ubVypblaLv
NWsMiJWUNq0HcZdeDfYMPjECh8OpC8S2nDTYKgUtH+Pi6wOkxVg4ZvD43EN/pirJM5rX9ZgZvmB8
TuFzJyl5JveF1CXqGKCxMTJ1E3SdL0u5mRDindgSAMqASfKmcOSEEb1L7Jd1Cl6NuQDmfuAeLMEW
xRCR3lOsgiMRSDrjQexzbuXiCjOXjX7/MEAUD6/3GCZCModjmZ/0fFSw50yGH2DPSEw4fvR+PaiU
bl7wWXcsq8zd7jwz9qBT2BIWBn02P7QGrMaJiB6dgBb/nVPL/Cs9CklIAc+klHfxaEcLUeZhduo5
9BiekHOMeY5aQSSRQyiCJfQhTq58jJUGj3MaqTsU5HEWQ48cs2fWpfHKAxFRm6wo70GxnwWAemJL
NwMC92rw8Z4DElkhNAejGSmAaWKABUTVtkievECRYYDW9o88YYBGvH1Xyg/PxMtOBaghHsk1zqwt
dMpe3W0ufZayjYLakdAbZc9y2/toXvT+Rynaaeah76FEy9yoWhAjEYbmYMb5nw7/6XOkupZzaWkV
j/kM79a5COVEKgCprtgVELgUEowGZp2ZK+/xtBEHZZvXVsi7wrrV0sweg0WDoyJJVf8wOWPbw3kv
ExKO/wcFJLA/0Ml24YJCUto55Wq4jdg/vokbKgVem9guPuQwL5KZSvjlcmZ/FCQ71z/K2sc6hoRI
24iidP/Q9MCs9ezyb5ZakIPp7CjonomKXLHNzfgEAAu5SdmP5/PfXuenjFgSHUruSxriSaxWt7c1
CMDBVnaZACEkHDm8OB+B75i/cf7CEc/joMwah4+WlGUbsvAhQ83hHiDHGNjQwAnbi2gHXakTPyC0
CtpxwXF30s7fGnwHnWxj7KhslSzPIkhhHiImqeDcRmPIjw1f87MKybkrpHNSrIYdSc0327k/1Kt+
pkv+lYmcNZ2CgXpYU7vEJP3+C22FtTX4ZSmWl1mfUw83fgjqpmYe82rXOsHgqs0yBXLErS6Q24TS
LQfYnMGleiF9+zIk1lR8Gd5OmdSuRkAPbe2uY37nx+/J8eTWEcbE/jqgVLdxPwBLb/OvdkHwEz/h
VxdsZrXYqUjXR+Kp2fnxnXgiZoa8RtKTYV1jiHniL4D3pKAth92gQcZoDA9WB77fv0GEVllvKNnh
mGcnVww+DTUWAyW98qoImNgZP+fTEXjNF0xPWt9yrfzAdPkjslZvTYcx3jJOJ4XP7vO1POfiDYJa
G4Cn0lalmgVLX6f5m0RC84xiISj2vMNbw2DxQ3huLq5GoOBKZvjbKIzAlLwc7vP+0+DegYGOJ7nF
B7EjK6h7K/h/YTCFBVotijFC5F0y+lsHxm6gDMUFiAAyTcRFNLX/vQ0tIsQ2LS/WjKSopoP9YxiD
0f+/B0GBhKg+k41Ecs+K2kEFHOYm9UQvkBT0Uytg6DmScn2zDtmg5lLKm92YQJ/fFjkLVERRmD/c
6NRwp1Ab58mfGgbNF52AdSFieAf3a02CpxFu0EPQoCtgScUrWiWhEkOfT24ykjoRnhkac3oH3x6c
AHb0tCvfQFq5X01kGvuLHbwqVtmniAHGjt6Vv454bugmn3WG+HrjK419GnsyKk5Rwl2PXd903JTM
9E+I1wHPylMLOjVDuFrqfW61i+lNPEG+Gj/vpSuACL1/57Q3mtA6ZySB0dwZ95+29CggV9dPrn8o
9NaaWdnuw3CYNdZk76nEZhxB6e9Rwtbcv5xUcyeJQNQm13heSLF+bVfknM6gyTrhVsetk4ThAjiF
hXmlppugEmaXlmsXt7LqyZYdr9nPu/S971oAtL8gH1yg3sgmJAddpe9BkG8f37EJECX7eToV5UCE
/uJi1nOsJRd+NbD4TKxIEHnHG2YwMlePuiT/5y/1L2hTlgf9RYSN2j2Y9nA+oUfJwNJiu7zdpyZp
5um97mS5lfdm3XVTqV/uFEJyOhGnpi8ETEETGKJ+m/cTVkoqkPBWQKzwGU3cUxR5sZ/uh/f2HbZT
80FJ2DhVEe3791JQL1no7KNxo8dyBFnswlhM7gJV2Vc/QxBJ6TJQSXzWjAuG66DNrlOWQEbMLF5E
FSTdEG+C4Uy+HdRV07HtPfFPF8YFg6Qd1dRZ2EZhHKlsRKFrsA33MKnlydSIl/Rc5zQpU0XVu6ft
9gF1GaEBAcAvqahzPQm6/3UbiSNAoRSvUpdKDHRSeoiNpwvCRJSwO0HQOISiNPU70G66QWJvJxet
mqYymh/9/o5Pr0sVilnaQeoyu65GTHjDx+lburXaJascfsQi792dwKBH4p/GP4uPmCFsZotEFtGw
X8pdfASIc70H4W/s2v5u0UMMLgboMnhZ8uUBUl72/ZQ7TRwFTFd2Sdi2f0cMQZvk3+8QHUjlwTWk
Y7ESwjUjiK/NFWNiB63M4aG6PrY0+vmU7esx1483Z5LPFU9GCU8u1eyJqEW/9KQ3MgdQV8BiTxAA
gG5ySJRahEJHNd1OB5RoMQpfb90SVsJ++miD6i9BBnQxV5tf1sTbAT+cKT3F4NWbgckaCuHpAxvI
aBelEhxj3Pmbg+HZt/CGlyKMfdjdNJQY3UjGimNHcdnzyrneR6R0ufGXwJzpSItjt29qYW8XWyaZ
FWSY6IGny+ftRSknSM0drkg15ECaF37PLpMHlCjA8CXxv0BvrcvbWsLXhV/peyJCFUjaGW00+AjV
Ft1OfiW0hu4l2Pkb4SFTDi/SdhKM9QsNBkHwOSSGfncxSjWSI5mrlk3lHUtH7yRVJ2p+wZtFu553
gfo3DTQQM+BvvaCg0Q2+SkG5fOPAbKJoiuyv0vWppztJxaO80GLEs1F4gPiYpz5gl+6JphH0W2QW
wm2WO25okdqBcqn0riKQSOGhZ+sc9Jb+0O3hi3pQ1r7IBgHRjU0eI60rv2q8ifi03/QvVO4lJPb6
BpwhHfWor+p1Q8KhJZnR2JXBrFvUup6dRx6sEckwEMYHDpLBCRWU1ANB/1jEw3mkvQLvUc38ZrDn
PtqLgbp/nq31tBi7AlYRb+9Pgf2v37ppqGNfbHaKYKa2frxNk2W2FknD+RWq9Fjd1gRa70qx3EQr
NQpXuQORUFmJqotLYe0hzXjfbOQfMNxLrc4aYT6aLXnZi9c2xkKAz0svzz4vaAUsqVppgO0cZ5Qk
luPjUhbExCDzpBHqBZ5YmLxWpOLfOQcipBZjroaLRsL2HB1NW00jtGuAeMGttvqGfxydaS4V7jmg
i1rdqEqqRnNNozwaTzzPDHy5mXtPHqomRPn93G9yGLO35IyDx4NdTycu5eYKt/p3F785LQnIICjg
eoIavtD+KyFgn43wnR+BrQ/ldAat3I7Kv/mhP1/dajB0X2XNKgfAcSYZeeJpMmmC+5GK+LMC+TKm
lOx9pHGbj+Zqw9C7NqPVhTeMtZN3psrLGdOSfVwvoDw4NMZzqqkCX8SkbXRg5aWJ1wpk/kniBpti
fIHIGMJlo1srm2pAyQd+DLQW1Yh8Ri4hrFZOiZpZSMZTjymmZQPvPGyKpNImrMp2v/LNV0C2Te3g
2QV9OpA/JUeAjCzycyKXHl+0DC7wqyEhiKm2Js0sEs+jf17O2Xc7mvhfjq7itwg5x1TmM1ynBR8C
sgUDUin4AWnJ0IIHmrYqh7jQM6R/usRvSZmrHOq01mIrUJaTtAwNeQTJtZvS69HheP9ASgbmj2Ef
aTZfxYqzkjXR2WJOJyc0cwgNb0ZycR/VRoUJf/iGrUZYEbPctqzkZHyc5O1aBXSQltdhw/X9mFng
yzu7yMwAvuB/sMW8lnrynXIo4aVYdW6L9WZq4JFwN7LEA0PYJX3ImLMvfBzKFsGlH8IJWhvWusuz
UPR/Sdt+TbxUOkk71TT6em+1VfRbOAqad48cX5WHvvoALdbyvvgVTM0Kkby/KcOalhCRxRUMUZwL
6Nj53LNh8zjz5G3oO/1GqHCe854TfZkmUe9OETRuUmm3aYjEs9gtcjK8fMQhZI19MY/hV3wk1tEQ
+Wr9/hE4cJIkhbStyRYhWz0w9eR0iJtRg6ZW6XVGJkGjlKaG6qAtbohKB0/zOkXKpgRiZk+Oj75B
r7EosAHHT6qYSh4tYXG4B9w/+di+04S+YfItts8dUqORupfylfNc/+8ywnMh59jimRcyuSOZ+VZI
UOAB9r0n0180W7CSZ7Jz6PV+q0o0iwdRS8uM9IqejWJOEL3veX8W8tPljC2S64F0EC/HlbMPzgjS
yk0QmwjeGWKHUFDXh52NVfdlXYp40ubTFitS+HDwfXViMdms9RLTOM27BYXJySViuYDxLB2wUM3E
ACW5s8KiC+5zUXiTchvpYKb0FEAz2RERt7LdoitOS7HeIRqPYaNvV9eLsYDXE47dazxTa4QadRAv
9C9GpbiUQR7ZpRQsGOPBsT1gLJuwR6KKR5nt9ffXkpLJ/hPa9R269RU3hi0DF2/c8pLUoLw1Jehi
S3/0SA1vscscpvy7YKeIc+5BnXbwBPPmCqdH3QGhyPVPcsVnOs30+jB4pkPxMM15Uc+gFudspBwu
RLFa2mtWhXlZjMIBVmolBp/Cu2YqRBjmtV/GIUmBd74Wbxazx2ee8QUJ1UFx6ugX1ayxUf8VugPJ
dDl5pS5e9k/HvO7Rk6p1u/mmrD9Vx9rhwyfYgfVeBJYZsFfoFwXhonyZJiJkRih8yPzkD+Qcos6S
WdjETjTiMxejEyS809Ks5aynsxjtPQidIwrF5ZNMUVe9L/MxwJCOoMGWunj09AOdh6OV4HzqR0Q3
ebvIR1xaZoP9dsy2OFDCD5a2DE8JPl04onAmKX16Tlukqw+ol3Qhbp+UAQfrTvYQdFXOAMi0blu6
8+cwa2wS3GmDx0V3vJDCf2CPIeNH96QunyDcOhrRKxTZUWFerw33mcpa2FCNL52A8rM1UOU01A1Y
kZQwpu56gBeM7t4PG6OzdO4A/albtMsR5Gng7oTaNAeTYTwHQpvYfrcf4RRovwy3GrJKXj4iGhMu
WFVdOITK2scD0Fh1dSMuy++t3Wj2Jhtt/+NDQZQeDcxpajx14uznAKRGOoONaT1QegFnqpvDlrsv
g86vGaJE5kvn4FwzSn3KJ96q9dOv1505W6pUjNpdJy/dTcm6yfJneashgPmO7v6MVmmsR1jSXq4h
cSGjIVnoA1KBbCqBWwmIPxZvT8TJMsymlxCmUCJ9y8ZQJdtWAeKspuOak0u99toKzEIZCI8siJTx
2MTT8sRqs6UxD3H63LKeZYe4RQl+9T1nZj1PMbZMYjUAXQQZUaLQuszSL9nzQHbsqtGwAuY2NMQ6
ODWkkizKH9Dh3CDRpmnyTX0uxiUV8QfVvGTtzQE5ApAEO04vTGlOaYsmhU9k1s9vofVQ79e3soOk
jVi52xVekYk3iJpepZHW909XE7qtauI7BKjTsAOEtFxV9xLoX/rDST0xVDoaagccbWm+FbAcGdA6
HHNgGWbNQbSJcFNaZSvYZdZfzCe9puNUiOr79HpCqUhS2V0+3Ojs+GUx53HUbvxgwZpQ/3jGBJPV
cMksEQembrqLzbVndlXbQkBOtXOR/WWBrdkGcGnuz9hYviFkiYH+6kbAII77QVgT5qRSr3WsvWeP
whudVDk/g7/BMmifGr9Bqt4tixsmMDLQoNj2RgdELTxguLSdXVYZpUdXf6/qn8oWpR18B/86h5p6
30Ebu66O1qCc1/Lskt/SilJxz4SSU4WGLFMDqbnZTMZcGZB9+jwJJXPsMT4WRIIpcVQXFdkJiFsW
Yp/A2Y2T2uwhjdGcOSSQQiIBA/OuuDubbkIF7C6mPOFjkrXCU5O/zK4QE6S4gIpESEAsSMxlZrpU
yT3+req7XIk243uEXSVpIpqWIl5iEeVAmeq5B+27rxkX8IOfoE/XCsTexXloV8KUNBj5nwDU+DBa
zCPHGqWErs1bNp0sSsESu0HQ0SNcb6F68dfZmad/eNkK8FQxuLiuXFHH7CQlw4RRPh5a5sImprbh
ErrHkJ1pPU+h5Ll6gDQ233ZhuJeSi32PZVcCXOAAx6cVAZ/4LFGUPOOC1ADf2NR9lFSpb9BsJRH0
/BxgB0KSLZN9zko1zzapmKs1siW8HWnGtwAfao8PHFDCa2CsDIT97gXaMsvlDTXYB27tYe/9uf5E
l19ShV+5RONMVLhGB8gM18Afr18vrg4pbVkA4R/HHiNNG/ealzs/sO1RhtO26JA1umljzNEoWGDE
PCUF4CQ+jrmNVHsDdipUzI23GmhkbYurHG47c6nJSxHEF0FgSu2qFMCwJVHsi1y5SHqsnngLauxd
qqL0xrK9kinJgy3nBbGKgwGIIwxsNDdEu9OBAO8cBy7YUFr2HjZp7By8ob0IMdgxGWY9A7zOvVyd
x0KL3exJIUbf7pruoyRdPD1YhpiF5vdjh/PiGutTibHHUGx1lg4+2Rkj4Hbbzem0/1m1yCvXIfT4
R0kGpk4y/2r5Wpx3FeA4RiLSEnpmeZyB5iEyigk8w6x2aQ039I/eVDW3QfntIgXFukHeJpOijD2J
wLg6SCozr/zo7vSbRUtdxfpudItL1rEDlhw2YxnxvHsu5Tds9+5g3qtKTjVErfdnf0YuA5uETNHK
gyQcECZGet45E5pJhE4bQLX7sF71neXu8wMiZp/I2avCm7hYuBqiAoOhtMMwGDnNURoeLm+/UN0k
0mmGvOT9AbS8XiXtekVJxyWKlRHLc35OYn+usnJOrDlTQAjg9nBQFOzPCkIypjt88gnGYlIpnLAV
bp1qrZiMTvLboZ34DrPszhK3sDEQt0b2wbFBZU3oQoz2guUaz+majiSjVVlBD6w09WIXOmBbWO5M
m+L4/lbNKUCpbDWYgWNpR4jvfF/WmmYmScFYbZGwpzGrlmDW67MS8pVeOvV0NzHGkzZP5RGRB56j
lljyA0/3RePsV9S/z4froQ2JaKU0UKwiq7zgB6+a3fjbYLjS8pH5Oskr0/cQNVlAn6KLCjfyCAUd
76oITOe4Gsn9S4U73qwG48mxFxafOBDle0KNeJIJUQWp41xwJpn3iMn8TsNBg28MxRFLbg1gP10U
GgSIR78LXsPlLXvuQ7iLeyjo3C6JLoAEHT0Za/hi86xru2Tpqx/0Y9TFyTms7635SUimgt4EemNH
1yLYdmd2tlYeQmOfpzWnGvsP8HLKGxpF9NwmwR2jLseZ1ISjXExlGxg8/5gddpSDUdfPqSjrasSj
1gotLMT8LeFu7iBfMMAmEzfbXlOAJAOQ6NRY12F2Q47Mf09e3CZ5Wk9ywpgdeOtN8lQREWQEfzkU
cYgFd10lOhTIJc6xGdCDyq8m8vWoobNRRw6oPgieyCkUFnNHDR8fOHtIyycKw0DIwrFYXFsUoos4
Wo8q5omN64Y6q1lA0K0gZfkD7e5C3+CG0PH3dByh/2dVxNcMqlqtJiTvY5pshCLQxCyZsscmB143
UkxIlMkEQOu8P368iMtWt2q6zviRCbM5hvLRMaLtnW1K1wow74zsWhB34vlNSE9L1NlnBUyk3n7q
YZbnrSiMpnfDcDkJdm3URvbOjUVs90Qcm8NB4/BfNzH+tL2SOKRcWy0karIO6N1QIC5tptlRfOQQ
5S+JjqqNZn/mhOslsiA5PEdus7tBNqwF77z7Lm0gFugLBMTyz2K4GoWhpbLym7wc4F6+Mc7pkIXF
Nu/ILYecWL+kReNEZPcMvhghmsr1MVGwPbl0svpM3UZrXaH97KZh2EdMkjFox/Dika+59Q5Uoupr
5X6MZ3yHdicxVunuN+QpWzwEc8kLCBxUnLZnCtQhyNh6LoqG3JBRUzIAX0ZTBLYcn+7tV7gXTMOP
0lE6J2k4rnTggD+NJ0ZFq4XEpvcpRphP0Amhh4OgD9gEFhMlYHiwEWzv0BjuCFN1ujDoU4LkRDPQ
Wh0O1myTfYvgNvRVslORwHGiumSE3kSSl5IYElTDk7NIPtaMgKT5V6FELCZYcpY39klC1v7P8FBD
WUXWRI4EpADXFyKr7s8NJIC+Pnk8t0MDUiX70ekxQVXxHpoVpe4ruCbuGEcpjTIx+LroWRBZtPo+
V53lrXPnXQ9vxuFQ0t84mSIj7T09x02IjhR/wx4ICTEJzJh8U/qUUJiHhWxpR4zRe4jkHEGyZE79
iLEdU4yKAjmaGL4EzyZwQfNiYpyRgEMN21/9NgW6sTkTQYgmmhvKgewKnGJJWH6zxZ9hePtDvgkJ
9r0neI/4cH/vgGjyaNB9z7uryQ8iBkDcCeNLQ4yRCvc4RbdgquITps8wLmJMFPwxSi6n/tTeb9Co
KvZd4N5qwe/8GSzsdiUB2G7OdtKV7gh5C0M/IXnKC9zFtozHofmeUUISXgjq39Hxfs29VGAnaH2Z
Aku5hoSuvLnKbldd4s22qSdgx6XTUecj/+GAOMg7trstrDD49F7yDT6IQ6YujE3hXTkpSQBiPcA3
XeeA8W3R73tiXMin46LtfMFEY9gnQmzKYa2omamE/VuGC2jMIA8s5NycIME8wOdrw2O3OqQET1/S
IMhYZKsw2DRp51fwXrc+azSqojn37q7/8F4zTu3zP4QS7bE6+6MJMWvqv2kd97+h1OJKj5UH0E6+
/6QxOj/RJPxJHOhhQe3qyLL/73DkQgctVpuGGdmQ/IV5Ad1VdrW/wZG5ITlRcRp9NfUf+3uHdvDx
rmogBiIpPe29OZeGUDfdE+QSPX+dr1CPfbaBZA6SPwYlmwBUFedBqgHVqXZ0AndgDdrc+c/8RgRX
kRCuQblStBwznweJrKxZ8zK/7mhTFX6WcuM1vKLQAxPvJSEegRAptZWmvffZEkUsx1OZVHAc00IQ
aO4LayFCim9QYHu0sxeGZzIPsQFMZERhsGbQOYZKIf3vrobzZbhFcEIkQIj3aasy6VqgI6XSEIV/
4GlrZw9allxygrHF/GteaOx+0fR+VM6zBhCPnctUGnK//CGCCgQMbU/zRyJaxEzqG/wuJMmcAHX8
sWpAZo1zi6Rr7qTvZA0stgfnnE0zxPek3UuNe2CN9/wIHBMkom1stRYsW2yVJToTaGC2u7MEZY0e
JYWRsJg01IUxdiEPYXucYaAh1GJ95LjQGbNHn1DKGVy/Wwerl8toJJ9X7okZZaH6OtUzpkPgDjiT
9vnJV74fQsXaizE7hcwdbpHZ3P6zJIxzyTpglRyAEIyYyOcVsFrt0v7NvXOm6qU8cq16bofHKcS2
n2B0RgZm9c4wMyzKKZSYhbO3z1aqt2bI+nvaSppoyyvsza1/JVAC9GXhT2nNPxT9hp4ocyYzTzZ0
NOJm140nx3ymFO9SjtL0HlLLs4j+dywyErjJFNlZ6CvDAP1XJkJjq6fPxDXOuSurW01KlC3kYK2V
bg1rJgn7CLfejdZaBQYZ5ZfM8tYw0MywtFpkLAj1+gUvlky+OPKVcRqZLdSjE0GR/1VLK9PA98v3
m8TdgWWm8O5+5KJ3Z2HBadMnVdKsI0LYoTAnzaRKltJwjaHzV/T6JMcoiSSJcHkXx7md/z7LScx6
PFTHPHJcHdsxDO1JZPMIn1PTF5WgvqAXL+1GrljIUje21u+7xrT4LmoFMNbTXDpS+5+mXWqfn0mD
W6DzYuk/aGjEPJrB3VcL95TUDS2yiGk9+Uv3+amWjhBa2js2ZeBKGpjWloZHLoTDvVilMqRncs/+
YIdrwXSJSjtLbJ1IkA0eAvYMHDU+DTbDcT/G7UWeXh+eMhlJ7gcRYn5gKWLEWPP6oDLBIBN5zbPX
NEjXMnJPRt+vCUDjFXf4TRsFqI2+YhI21V4vWevicBKhezIbs1qqhHx40/IpbZz08BzYkszAIrFZ
IDuJeHUD811P/OETGlNzpRWzdtOuz3+ue1esNfEOwx5FHEPfSNr8pB3KOw2Yl0xYHBv40m+C54cT
xHy2+PEpzYJh4JfnzWcYIGnfZp26qHCny59PsdVdeXrPQFkcnnad960/Ib1Vt97QyP1GVY1m2vMl
JeWm/I/U5qv4x4LiLWFhw6TCeRBwLm1KrRmhlGkNsHWUqc73PlwkSfNpiwQycMk6It/IfeVD9ziB
H/GqY7oeQ8esbmYSw6D6hJBe4ClHOZ1uAPqhIxijGayuym5nBljKG7GYXq7o7x16kU/2QlzZKrBN
ugFxc75TMr6kCYYLlrTmgkeYdNfbKIHi/DSAfzqj7tKnvFJcd6t0Yc1r8EUY64UWl38XZ3bBlWg0
Ckuy5F9CUWCl9GY3n6h/+co+CkqOJkPSWovFD0OcYbCQBue2V5g2tHlN/itv8SY7/vKrg23FLz6u
jMzAnT0WrcGxmjiMZOfZNX9Co4lXN0Iddq5vPTbqsIOuXEOfzm7+v05XCP4bWCyaCEDiN2Y6dDA6
m6Ddxuc1gMmEygPqkiNlNghex6ic9x+lfBHJACQXqjFiLz4nlnSrWX+s/29IVKtvuGLsnmZ47xXP
kc6rndOaoMaTYpoeD5QkcXDm/LULK42pKJ5Si3pqo8Rp+9peeOywMhQHLAkXQFCG34x3wi+b+H5d
pKYIMGj0a6VOacP1O26E5iOGe3R/MBrBQcD0OTgxjyL8Y6YaNvt5TtCZrsGVCm+B+k0CjY+0l+FB
QsSbeFs0BOnxvcOVKu/39AWz99diJt/BMbTf0iU0gY53O6CSZnWPN86W+R2xgVGLB45mmpwCaudp
QOPtuCIh6CxGomK23H21i2P761ZTjaE+tMXoV3OkEPRiPLdls+RaFj6udv2AuNcUqrNIPvSmr+HB
ReCgr5eNsdDsbEVVwIGT9TXMIM2paQ0fM3ns2ZIwP+sRdH5ivehvWEnWp1bNDIC29ZYaDQty3v2h
a3tGt5BYjlKxzJMoVxjGK7H/zPkoh0A+K6wyiMHW6zkaeJ4utieIMaA/4eZuTl2AnS/MyYKpRB3v
oArktvMrag8zxRYIM51hZYmYacBgK6ZkyRLf/2d0w/gFm+yjRQvm05Log+HOGANQmm/KbStBue5m
2et3fE4G3MZ/GSrsUX0X+ISgSJVspJy/nP4wyVtKapbyBVHOgv0BsEAuhKcyk75AF0+7VjmNZgty
1EYjph+n67u/HcZxKuIfJxtNtjOtPA2RGh9aBVkE9MXldvJCSDIiF0Q1vuE6UCvTXB86d0o/QBWi
hChCRe+ef3PWg+2QMzz1s2DnEz5o6jUXU9j5pzdjAQOJmnFHdRU8JDNSnGr7E2951nItFsNOCcDk
2RAr1cZlcaE/zaar8wiqXKR1E4vGY7WAqC0xa3cBP9Q2vSeHsFVfq5R0LdH6CkruWF8+SLBXASIj
B+DWAOyKS/hoBGYqpa22zLMVmXwTDh5adLDCqb87VcG6tSoAX3CAvkQfahYv6yYOxfNsqPNwph8g
QleraMHOg0hjQrBZxOZzs5jow3YBam+Vev0cjUCtGr9KIezGbkiwdUS9BNBsdyRN/keZwhZbnSJ0
09/uwJDrGXXaO0unKVFJlMWpYoL8izbVzUpNvFsATW4ls6+owL3JNA8DCDO18tJYSIuqUfP2mzXP
DmmMQDlGd13oKupf+TybEWPoldPIUIh9KWtIky9V6wyIPKrbXajMtHeHyNFk/SHvOIi2JEtEv+Ge
DmOOGgqXlr4py8lumpntGv8oSIETZPap80tIVFKrzsGr/5Uh89d4f1kLdPNKc+Ou9I4mnHQA56Gg
5MqpMzWzIjg/L+c9CNrmfj20SbsSrLuduIgo28q8yiJWb2t/JAbGvruW0f4G2HVL6fwSh3Es1d9J
aMz5N4q0FhPbwvImnAYqeY/TD6AEg4zDlfjMl3B9n7iZ64kBwd30t+1A2L388wuTNpjt0PFFnlk+
MFttx1mU3Ler5VJYKQL1WyqA9+MnrESZpQE+hMenYt6WFzFWymaB70NKTUOSB48rXnDuXUu6OGIF
dyVxTOtUWfpvHpf6rlWxDlg/kXHcQpCuaptko8mL1vy7eK5eItP12132yfQSV2kStrGPOsZOnP3A
4IXdZ9DKcJDHDr1yTxVhI8Q6z6eMag3G7j/LzdYAimvOGbi/igE21A4b8b69ZuFMTrFDxT+WdNhS
wHkLyERl4RkhQOHlcXZAJQzwI1PWQFOxuCgAkquBNA9mTR9Q2TF6IX22qFpghU8UGRnb2slvqaHl
/BdAa5Kpo0MTptD6HAsWFHXcvIstd3RjPvd+lqbICvxuhwXc1ZqA/8r/dCW8m75PQ40Owbmh7tQM
7yNuVU0oS3iUJ2zoHG/wzA3iefPP51rKd72KDFN6qZIqQ4ePPa0jaFt6oso7t7yQKQJzUAxcKq27
Er/vau7vo6xMI7BVH1OJcB78vlmnoVfW+BDrt/xYB/1Bfutw6lANYQ52XYzzxesd+c9qRaGIJVzv
R5uG9OQGSj3viU3sGGV7zUaeGg0t638FXV7vnARFdVzP/eezaU7LgNpWUl/ZUiIfZn33rLOAYtb3
2B1nsaleFuqndCm3ICykxeKXOB1kfco5/J9RV4jEYxfu70edHV0x4+sDDL3oQJ8xGHnsNrvWh7dP
F8HwFohcp5beebNAOaFiUlYgLuVSp3yr9xD3nFQ92yWi0G9lYLfvRe+aQ7Mry6kxVVn/s1VCcj6i
nfS7tsBstTMK3VlHYN/dNi5PHu+jrBDp2PMdPoxVrJPaAGA5cvxe7u3+QxK7/JwhHBLToHhJOETL
l0pCgVVl+YuLNBqSJq1CbJjocJZOqyUeBYzSokD9cA5f7uoNtZAzN+ICTY33OU+COv5Vt75FNpFK
UEC06ihv2t08Aw5TYpcZSgxjQ0nQ5X8MCjD5nNblx6aHx1/pV6yWaig4hzHaoE+BjO/eX9o+1lbd
U8ZHhLPlUBb1Yl6vA9yvvbBSrdM8da0YGk/Jt7qUXRfCWjO82n1VIQLhIiHal7SMnRcAhgHitXTp
X9tbHJKI327Y5PSN8Fy+m7I7HtRsBYP/wcmVYIGnfHmPd5elDnzXJB0HsiRCSh4t6UtqN3CxQqbd
LviY0N366dfWuh770yU6Wj2l1H6oR1XPOqoAbu2rUMMr0vF4hFl7eM3Iqkds/hS/Sx8tJ/n92EfD
NZSz9LKvDCrxrKVB55lktbqAd07h/PtRnhdUWWE791InHVI2ztx82e6JXlrCU31ITClKwub8jbwU
wp65CdQOJWRfsFXwHWhdivrJnRImJmjuNEwQex/q5ei3/mLT849XMThL7g92P6NvRr7OZIEYQGsC
YYy2uik9lcXfoV4UK/jhtPVnhTRGEgJzRuo9ZvgSdRlx6tt33BfAptL37xMu9OiKtv5AgHuSKy3k
27eYGaFwaiiFRjf7vXvJPgLwOVaemwjkfuU6/15ai8oNRlwpHZ7Np7O87ylXNPoBFqG52ZN65Xu7
qtsuMdRM2cUR8XSlaWLWUj3v0w3LEo+M7vsJGqSVSc2LfjfeTOZmK63dCIR1JXgVqNpsCcLwWzuL
eDazD9MHiaiM0Jg31CNLT6VnHtUkIf7yaeWHGEa56HdcxVXCBzt3th9glvg3AibgdOhjwg+HPRb8
Dx3VcIcKCjO0C9U2rjB0DfeXdHlSPAC8HSrmeaqRYtiz3dkOSw9hpQEL43xmlxW+FYWy3+hrxccK
amb93XeCLXIHJuvAS9zSERKBTXm0xJmwON9w9ItH0+C/EcC9T3nJh6HkLZtvVPUWrroSRND4QwqJ
VrD1+gEum1MxjB1LlW26itZrsa8nc/Cvv3A1AzEn5JfGEZ7shq8HSlstz/Xss4SI7vCflC+Os9UQ
+S8foAPZplRk+aEzKr3UZnPlUl+Un3IHyAJRMyt8rrXjOyrfK7Ojt2nZzWFXM34RlOLFR6zmn2B8
K3hG9qiqmRh29tjbD3lwuMJBuOdMcQUvjyAsV4yiERmLxsR+Z8zfk3fgzAcbshavqll456iyVNwy
fVbKzTPvfMpa6cQWiNyK0SsNGJCGwWPuseb5jn9eElBcnr6LRhyBTfoPJz07KTMatqOYYmRmSQTy
Qmz7Dr4RDSBtXAd3zT/P0kLZB9Fae6Bw+5LxxjsLrsZIftMxlhlsMUfLWRkOVAiJNlaJnBiM2tMn
Ke7/11rfGgt6eyeXhO6/7PZO3OqV/MtHFPv6VgwDjLJvmluJ5/AYuU+RKhMg7jQM/p7PS37OBeUJ
vnvnR1NKhZpAfwNuUMT+oIlk6irNhnr3L/m2LmlsuaUqc5lY3FkEWjTYrZ93UX9tRCf2aM+Nywgk
tF2B/Jz361drdCs2gUq5alxsAYwAqUF4CbOjm3o/XdLH/lDVS5mNSDxyoiXMC7Oendl4/cpo/Ae+
y4kznktG/+HLFR6vSdfSALzB6zqF7jC1L37MAIECEg6VB/UsLtA8FeHfN2HqDgEp9R2oLV6KcuBd
v94XcoKrGVNsnDWx4P1aE5gBUyRjyliJwWbtqVbgIibVb+rqXvSzNQFOmjY5Ac72SLtzFI6kyDGB
9dR1KXAkEjc/UX+TT629iOX8U74cpgsl9zZGhYAmsbkI4Syy/tCb94Wd+aWB2+gfvtLDw873F47T
vYudSF7enVU05b5hVrxzuJqzGVIwxzw0xnUC9WN+ND/V2KPjTyh2cUFH0lwSG1WZjiSVAFyB2Aal
FaBfTwthsS/oWKVeo+j5UtUzLdfWQ2qvkhGsghH5HedH57PW/8nJzc36rt5J6QkmrffQ7U5EYE+H
d/29Q/d8ZaoKDfmHd9H0JsafDB8WxkS1sGpE0RwSao24v4uKE/v8pGkh0c34OfzSm2Zcsx1y/QF1
Ea9ddseGgvvVeLna9Tg1dNWxDE7C1FemTPcO3Zyxh7MvMMMHKunnthH75TMUctzKa/IHKfeRRGzO
oVMXals0GEWRL+/YTEUo8iJPMD3iN4Oh5o2W6UNuFUN1+jP9+Tv9CV5E9VCt78RbNcVC+SKX5n//
5iN07ANKQIzDndVR9uBcs0pbuuHTY4tLD7o9e8XY1ELDzrQQj7gRIYXpKbmEw7bJrC6Hw0ag/DUa
F3pXrhCvJlG9AVtJ0/I2liuE6J9s1wTS0tv8JTQx2kdrT9O0795hCiLjJOvouJIdNY+1d0Xar8Sc
hlhBZsXkTZtwnBFVyaaDgwJVbcK6KxjRevNNBvkOZ4syrfPi6VIEwE1CvpWHBZcGc05TbZGK7nAy
/JshzeIvpzopIbJJAQsEKFMYEpqhDa9VGdLM13gbAfI3Sg38OhMvuDLWMeefqTggE2gXlbgqgSkz
k7DykDc5MvWY2JoKAwtja7+8lP53b6h48uKQB0OF02FhaE73TNQXZQq7ORQ8Qbqlg0q3z2mGTLR0
JZC+HeJvrleHqRk+Mvh5fXmGpCBNNVFPbA3IgxlSwEfWa94/8s+3bb2QtwMLEkB3qqNsYJEvRphY
Avvhx0UYQHrTMxV2EJ/58i3EbWuVLhR8lwK6dfIewE98iCfJtrRfk26n81qDUG8tvepIbHwjb2sj
2HyigdhA1n1mX4OLVtNSQref1hytHdcg6+XP88+US9yB4AcCqUDZ7E5rjXAgiay+h00Me1RGlb46
jqD/6p5UDW7S/rHGA+aM2Ll8jr9d+aC1ukoonyeX9NC183zpKLXUw/DUW4HE/KOuXy8hOcRCAlZu
8bpN9iyXcIpEVUTOsX47vL4akLSTTKUbq8Zjw5cA2EIk+cmWJP24L7Wy6TZhAti3TBP94AHrnOlq
1ZX7cJ88E/l3IMCqSw5fUATUYfeiGsnEeBLnTg+jFkMKGLJuHyk4MvN6Es7O30w5FJGFx9FKir3w
77QYGa5VszEZPeQO41lMOYfkwM3luZtE0mO6FMFm/DQVyKvu3IvP5cY7NjrJTXHL57D1Un3krqIG
E9IWeOKuc4m/L5E1FyBLDDwymdfPnbutcBJvHbHC6tj+227gDNTpurzE3pvM0f35kvn9dX6+a72A
Dkx+M/iUEjYdj9bCBUIzhw7GK4izOVf5C0yoLxvc9n9ODqIhV9/JX+RkexO2xKnzho2g6Caq13pv
lz9wvV2J5Qii0yhX/hfV7HfOw1aFNVI9mHAL2DkDNaZn9ZC7qBhQfDGNmUS1vHY9H7x5F8eFRYkP
e+/zblGTT1D8bGqWxmYMhVvetHHC/MZCE4aNTYPCEyXYIbvEL3XPcdSQ9mDIiQau8BdMKQ/GIPiv
5nahkHw5f5lfE4OUHURccV8b4F3yWwMQL0JJHwJogS5DGzsUN7weC7p7DCNBtuzpH7Ujb5B1rpXB
PTh9MjzWylKG+MT858OboGAbEy9GlVqajwqlToco/2hYIKQfTnnUButXg5SNX7izdzdMzrxvTiq2
GHVtZWSuCVWWfPYfHivAyXva2LmUe96/ZwUdEXC59I4BzcuBsq5vdMiwv24eYwfvcR4DfqVhy2YT
sIBvZDuxZUE2TWgdxUvMyC7Qu+Z4X06W3r8Z0BN1aXM5pq3Xizx6F7JsZjXtaOSBpUqFNFLTUzX3
5tXu8Eh66WdByj1PhlREWkOI5E3ZPWz9pKHy+/2GhbaG2AuwuVEZ3f1CZ780/c8ag/VoePQTmkYO
5dxpdxUxRV5s8g+imchbUkmtr5C5okFeBxo/bMVzjI1gcPygY9DyXsk0f46nkZoNXqQ7DUqc0Hov
euoqPpobnc5xAcYJ9Jek/HGf15FYBZ/tvogsgG8lEioPQCjRJG+VugdLwCx2mj9csjN+EFpr9Mm5
yvyL4Kj8eGYVr1j3ZmVKWTSOZSED3tIsNeCTAkTB4TVuYzkr3XYBNMuyHGG0iRI0zfos+QB6S9MN
76rjvvP960qWv7IgwgDttk7w7xhO19zJV9am7KBWKJVaAp0PtD5MT/I/9Fw2Hk4dCS3xXWo5IScX
H9zk+VUnuvUUDZDugXwxREUVEhJt5se0pUFXSrC8uwmaE3YxIzDe/kHERdWoS36aTQIc4sWvP0Qr
FbNUHMkb6Hq+prjdr29UMQX+Ts4w8dTACoyJ2h2O535E6aOrs+pYkFyqDE3ZucKU8PsyhiYZgVfw
veFelH42WyAhbjR8oTmbf7CzUs9OCbaGV3CZDB2O7Jnnz3Rc1Srdi6xi271giWXTN2DfUR/QMqgp
W3Rxv+yBB22sLXFaPkWgUQLq+mEItFe42HNddbkSkw3LkZ4BOLQwikyPdOTno74xFmehQW56y8Xu
PD/VOK/4RijCLQJVFNdHhFd4p8S+fyAFhsYzR1FzMLeRrhawEcG+LVqQ6iHZYX0qhYAmYj5cdLVR
I4x1D51Xmr3y85o6BDBOcDwxDv2a4pd7Mi03kPmw37SfxqsvTxgEvXO2g/jqlmwdwh1g9dFgrqlC
hoiN4oHDgIPu2sCdbvOs0qPCU07UeTcyLm7AwaTKYQ+4WEk/BddFZyPIAEF4sAaXx2EYWOhocBLO
lgPj37TOrbEFufU8yyvRkb+2UgL2KxxVoRJGBofJr0fk/NEe437j1RTtOcFKVDXEp26n9vwV9ZdD
Oo7herkKP9+I8ADaMFlkvW4xxbt+ItrJaAxpn0ckwhLU6EOAd09nqTH2WGlxfMWhNfvmxI0CRH6l
sUpnuMobdntblT34aBhnYkKrhCgdXhKquWfMbTyL5RRDCSH3y0xAu6I/vYfeZDybTAv3PlR4Gcds
hyq/QQ/fKDbObRBE95V0j/kLqxQ89n2zx9mSJZsde4k6s1+YPgIXHVNJQ6qdzbV+PWTA1yZ943qm
bfrr2PigSSQS3MbnG6zdyBCarB4UD7ig06N1G0vXecYXitpLFGKWGxna4H72q86lL21VN//aRnIr
1Y2L99eIS0S6Bt/VFnUAOvG90DEWtN5YUcTtv+KXQBHImaoP1nQSnHpl+68TrmMI2QKan0qTQe4s
6Vik/Q0wx6dM/ZCWnLg8ODIh1rzUnPX35oxiDcCXsq41cgDRDJKte7IQQ2VJ8s9L1jDRuzi6yYD/
oR4Cx42Qcuh5mQhrJD2MEwz5ifEElT9UXES5FYndMziYDutpNKKXqv1f44v8KLoD/E0seDERZHYx
RfydSZOvgzz0/pnuOMximo3aJTJjMaSNZxofS2hWKm18sG0s/uaJwFLFYR/Kn18dx81iccLTnfOB
/u2SyTBreQxH3S86bMgpFONSuRuj779Wiobs8o19w7Z/QzvWiwF38dMbfrs9KtTrXfduiNrt6rzH
WOIDWzOQz+pNGsgCIfZ5u7sHRv7MESttq6tqnZDJalp0rRTNkg9ucZsBtince4ixOm5EosOnnIkC
KoyeXZglRkRJlZ4W61ucjFJC7SqC4DRUGpCAxRabk9NC2IK65Tvtm0mF1REmkjiecju2iCs9hjWn
Og3RpQdNWCTM5LO4n4Y9JSZwHd2BzZmiJvxWOdphlMrZEJURx69lbhLiJpjYFD0K12hWoS4YfI+3
y5xNAZ2fbdHyZ7ob/f24tfNdTBL5WZKX9NhMdkGUZTTMkf9kNGi90uHF9XC+EyXCzcfzqgAGhBqU
Wpg6vhuj+l4TNthSkmAsTBSHvceGtV2VVQMNKt0wuA0qHeNGkltDh6v1MOgzADiw0JWq2qHIVlMg
IiFDP40ntvnSq9pSf5gjRmmS0n2LBYUeB2u2BW8zOI2i11mUtagduXvs9F/TWHl45K6Oz2R2Wm3d
CoYwCn4dYGRRwAzfXoCOiPy2KVMqrNxRanrrZpeQH03hqQ8xm6FyVAJ3OahIY+0F6P7S/k1sBFem
DICucWhOYPV/mRsAXC0vGI7ealXRIp5/KAUdkfSfnPkaSyX/CiPvztCwHma2FtjqJwR9BMzlYs+8
qYmkhFLhgWemgvGJXkfMPc6+zr7hx8Cg5PckJ1l83Zhym9QfoSluFs5lwISkSU3cNRDsYVpChdbB
DAek2zjDr4VPR90TVKSsyVc3TTO5Enx5D+E6kI5T0BVNo/A0W+enXyOX12YiyU1e9UrkyCh6TICp
jNhAW/Kr8vM8SRqoZFW1B3qIAo2k10e8J4PhDVrnWHw4+MS8ia6Av96+T5DcfWsqo2ehrwHnS1RQ
Kto+FqoOsxa+CITvXtwm7EI67jiFLpI5/6AvMq9Yqk7nzt4G0dRg/eH6nu4TlhkT69x3l3Jbojrl
f0H5w9VbFTeLTptu6rDoSsCR1I9LMgVa2o32Sr8ti7WfnE3+k0dyT1G1RMiRRWXIpN5/+FcPOx13
078Kf9dZ1Hc1Dx3AiocELBsO9oA59GETN9tkKAeM+0F1EgH/hNSJzNPKAmx0l9DZvoUUHsQltHrD
YGyuEddTpVseVlXx2K8fYeOG0iuA9qUXxX+LgfWsvoCsXqAkMAJ5CuAGGQYi9IpN9qDLHQp5vXMV
NBNDA+fs0onW+GsKUwFe6CoTdmgWx04nV5CvSR6r60ZNLZ3anwoOHdBD4BlgnKvlO8W3J0Kpgx8K
2RzBmjOz7DuQXW4EnLEnEsaBrpK2SaXCcfDrIxPxNeppd15YPI+IRCElJLkrpJX7KWwncKNIjJwh
vBL3gwdJ9nP2zvNgqq/R/HYmlBpd8FyMTDF7ia4tIYs9XyLql4LKDBsPCyezP6LDRnR9nh5tSuoh
4zjWLY39IS1kPrlztq6/kjxO035aX6c8+GX56gl74JQiIJKV+ZciGjrJmdH9P1XEqRsOpFINbCaF
KgZRYQtdVqUPQYXQCR7UNiEsjOdKSRoL0y8P2Ir1eYV26Z3hCda6O8xEcaUjchINEVKjGQnStRU+
q4T6oqUyJQA96miJgtAdYKrYp2bKjJ8q6WSHg/1AR+q4eeBStD0Puzrz100olY/Od80npuXlXAAC
BG51l7WNY6F65mbSghbOCfozojRQFMlYbdX88SyLF+YKgKArSGFbWMLDF7GThXZ6BWSwS//8211d
69BBuRDPdRG83qX2g8GBy0O/ZLFOoy4IfnsxHsfcwyEV8xat/Dm6nv9hXTxENJ9Oy6w1BfP5h6fE
ptJEb/5619o6iAaVL9UxxdiggTnN/k2ExI522rlgTtfKDSag5mAp+6a1KUh9dGpU6+0J5U1P2PJE
UEqL1UsaEHG7s5vBIYwFECyxtlokscDjLrCp3QLuHf+i2afDMz/3tXvNDVx8Qm1/WFCuc3XiU1J2
pPLHwPCsR44Nxav1yTq++a8F9Gsk6LHXVopXLkZn6dvg2BarpwLvPj1oVUwaBZvXKjw/XQBWyoTk
qBuMIMkjBq8HmCaNpwDRJVj37nMjE5j3nmFDZ7aLJzKHhhp8oO8Cj6xuwIHO8gLbpX+RDaUO5kK9
ESnOXFW5owX5kdHDjs4WNwahSQIxihLmzJy5g/OXHU9Hj8zbHYuz8kTTTjj1BPpMVnA9OzrgxYQS
haKhMuSagojnAZkVCLLTAAf7oeQT7F7A4tfPC+ncERt4KhI27rXmC/AMVfknbmL5AzWvmQR4H8Z+
x2j+foePjGSRMH4M9q79dH4fABkihwKMEeZnuMl9x83JOVOoRJxzQ8XJW5I0M2b8YAyXFWzIVK9b
L6lIv8CO6qysx3zfjJ58yvDO9pBam7e0id6rFvo9ZAZt1mjUthwXXJSr31PdE74dZDp+Xp30GNHg
abHniLCPEoLjVLI5BNB7B8LD6xfGj/YXpfz2ABnECwdcb7gYoav7jMDtaGvT9zDfTKby7bH89Z+v
0yUdeI0QcyBH/dLKVFCIddCSzgeiKk7v6baHrPe990PpAJvRVGHE9yBNEVLthkF4X2IHkg1l1+I8
a4JGdLC9d40Lk53NEPOChLy3WNxZDmJc1ooWSp2E+MhE6hHk1s1V1QNNv5j6uo15wA0LheLJNO1a
K5JetZoMxGeE9xDdnxk1R3lk+XepJbvY2FCXTebjV3AkoNF27Yu/hSFOZQCWHCZ4Q7ct7KY4yNQg
ciPqrHiTaZ/8M1Y61XmILn3m/IT1oBcdqORBwHHaJ+0qJEN/q4dob37PoygczASl07uPcz2pzY39
32vX3s+KQk97TT6I+KdqPMkfwElHRO9iFqyqSR2lYE+/P5HVFJZix0cptVs2cJK+STsGP+VZr45Y
fe/CvuHhl+aJ8HSG59oiqSFqvG8EMotIaDyWBiVZIDtNUNU6XyY4UMNAr4rt0aT6fA+qQKwb79jJ
7R4RX1igYxBVL3sKqqpWlNQ9nQF5TWLdD7GqgLfHkcho8MqzOsa0j+mXLfjjFu+gTsv3sWVs2gVS
C4ES+m22/xrZ/sz5ddmlbSbvaxGr8SK/g86tWTvS3Mr+ryuiSia6lbo4d7d5gstkbb0NKA5p9Bt1
iPxqNn05qCuDVIol3yxpY9Wzbmy5KSDNqx8UmkvpvOISQ+F+mNs6mAGy7+DjoZLnWLZCvXiZLfga
7qBD83lD4aaMgb3DnizE6+Tsm4jDqGlLTmP2xe8/qeogpUQC36TXx5oqk9w+jFR1NVASomfSO535
jvkBSkGT3/WzUhbqEopHFzLkrU/pQoz6fl2pBBz+VNjS0OD5Ukg4jgRwUdQiexmZ3JZXl6WXy3qb
4I2YWrIuaWwnuc8NC0w7QERDEJ9hWMiunlMTVvFrKEdrUxhgfe4YegrRypy+8+GnHXxh6+ZwU198
8EDXaoBgynlIbTT0RJNVuPBpQRxxE9BbkXnB+yf5UEBPoqwr5he1Yxh5uJHHqlY/sYa1PfuwiIkR
bdpillunFTiZ3GgtqhCj2WOQIRdgPW1aqiLu8BMDOWQBo5KLpByyHrtne8fgp2gzNaYuHoMzSTDv
ZlIVbO2ySWSQk5xLAKgmhtvC/Rbyp4T74q19+eGIY4vhNYdaYRLT7fJz2Fq746tXGRPSdAH0Paju
ssDLdvIt7Ptepq6q8+RLbSzvxpe8u25zVxJfqe1OLhYT028WxV9C+gietsrdfUCVI6h0fChkyoUv
d2gk9NOrNSnr+wMlDy5NiuxmF6DiuJxP2dcRbURFCWKDe8I7J6QXqXU8SsDlUP/6ojUYa8aEQDVd
QRwoKXGtQQZXXAVjQ9jPRKTlnLCfihBInsbptUOpnVVRKcYj9K160nEU0o2szjLlmZppaPKKlSXz
mCg3V/R2knONUIu9PMPJmXq7EjlkTY4NXSjlINls6745jB5+o6z+yKGxGEmv4/ypNMmrZwjlQtCg
mEaAn6pSiw0+ad6QZ7Czui2CSXYjxcRuGxwT4Yi4WH/c3cNgLBesYU9hNyJQuEkVh+/QKO/l01C2
ZniRtuyI82cq787oa6khcyLcDE5Jkd1C15p9qUTTzlMHcMvZYrmCl6pOowdpnVpCuueuWBtsqmSS
QpC/mYeiby3KPTvs8zK6zltZ2V4+dbKEWGlQoo5GW5jj/hgo8qrsSgzQZ2w4z88X7nWseNBKcZwn
BRqunQ1orD3MlFwZIjXMOLS8ogFPfCH1Qr4Y5gmBLlNohgGZM/axzisN2FBk64UqcpuVcOfyp0ZM
at7sgnIIoH64pH53p0FGP6AKQ/SX9ZIbQwjZi86JvuWserVqcFua6IdjytO4ZDWR7Ai8s2xidnOz
ZqmSFt5CS+3QttZJo9DNAuInP4IE7L4hTEtrGGBS3SmtPHah34UH1lbfDssKiqCku1/BtGHZB1nJ
dJGBltzXCOYaLZz1IRrxslEDjx7c6PSAJYjlFN3Zbc4ib6ld+f+ooCqO9EjKEEBMXXDWn7HQXrTa
zhJFbvzhOFGg8wOez6BJpWwjZl5ZK4+b284lC2GI2N0JQL46CNAGULwg5bGaqTABR+NecSYiyQFQ
S38Jp717VQbhC3IiYn61OHoTAhn7F+0cx9GrwfFw+TSBpDCXGm1ZRhRfSwpnalHNPYLomUQFswWh
S58qMpjYHZeEMwtPrmJrMP8IdRj13Zq5ZtkzHGXERY62hGJf+h0XBIJ9Udm9sGHoDF0M8jPw3Tpj
XPpheYYOuPscKLxKzgcmdRZGTHcooIkyVfS1to/MCdp8aBJTdFjQ2+UYAqwJqfSOT4/Sh73y7Uzc
5DW8ogiJaI/3V1/RpBrSq0gEsOxyUpcAgF8mrgSbHXYYmFynUw8fFAaCGidejSCX/lBDL21kWLyj
3IVj82/hT8DvO0OQCE4GPRZAehjx69cFJHA7t792/AuwW3AUipnIJRtBoTugYiYsmXfx8ITT9ypl
sbsohwUxvdUmhRtW3Y5xlHB2+7vVawqIhkFxtLaSXQtteVk/hwxTbBOzSIjUpqBAa96+mGDy09oG
rtsm1xqmiX2kLpMavMUTZer2bTEL95Xm57UUBOBunHMx/uoXRw8V6C3xcIpg24ocIn56cAMhLV5v
rKYbabqzsz/LKL36bJbmi7T1C01wWFmDje3IhwaCpXT6YvbDTlRwQoGscLdACeShvs3wnWD7e02G
JpGfWP3p8SjHRO/riP2sYfLOYqBMBxFJAMBuWwwPE0plz++7yzG7M67cj/UeB5XNoARGDu/pSvvi
JeErC9Imeg3jnQPl1/6Yf+gH76ZAWvNPVFOGZz4hYvbe5T5r59Ui3Rk9VTFoQD0X5XrNWSRpKIHJ
Zv/0CUaGtNjhDqm47oeMsjcyPmq1fSRwejD6+Now6ztE53O+49QL9/+PwO6aSoFnzMngXtOQ2ev+
Vb/D2nGO+XeQ+IjX/pdTkdmz66h5khMThOsySjf9buuFZRzQ05Fy/oJXMqChc2/qFGS84u8L5MxT
F3yHN+33Jg30s0par1uplTzDxDLOcV1gpXjq/4kvrB3LxtS142qPxdlun5Ug1AHmnERZlJ5t49V3
Ktmzfz8Km0Nqt1uMC3+fxk7TL6CPsXODXeS3y6LlmmQmfSTHQLHZIzUU3zsviBjSZrkFVDlfYZ8G
qWxBl1jtQf0s2qUNq6NGOfTdaW6byrhuKfBfaA9nn/LJksm3F7m8hNxY2l9IPFkTPj6kIL0KSh27
J6BQ/P+WVbx57eeWB3U4vTviVt+Mp6D4lUJm7jepjyBOft/F0c3/e8Bn5ezkB+lvORc6FJ0mkhwA
et+WG3cjWVSU3GBGoZkvEsx0Ss4uigBgn6Zafq5sjaYIuuf4iId9c84bptlICauW36vdGkk2t1Zg
oS0pOwpTalunf4tGO8hxXT3U74hpTNuDJj8XPkYd40inlXqzo0++MBsFxlGe+x1iD8MwooA93dIY
jeyXL5ycixwfbhC/ZKfFRd1mUzhFBlcNy9m21rb5WpXnW7SjHSaXPzMaKiLDfkkyLwFKWM3K7ZtW
H8ZydLvF3tFlNr9p4wrX4mL58vykUHi66rMrFiT/qrM78I00t676D5ZhzM2cQQnoYPLd4s8hiJqP
1gOJO07malJmt0HOItmFq7QxzwAwm7tqqShFGuYxReemwxNTi54/oILK1ZJSi7HCF1Wzrp3z7bQB
WzdgWUdqlpSXipm6XZ4Gcx383r66R17J7+cUfHnu2ZkIJSZW0MIizAUiVGUFbEtqXZqjmjCgCC0u
7wVAgmyw1GxOvOxWaQY9jczghpBF/LmmJc1FZ89x51YHGlFMWU+xaBrlVIrLoIAe8mh3CqaE8NnS
ou0n9RA3mKQERpglOXdKV9c6UweHH9PufciEvDl6boPgPTs0R7WMmd5l02W0rriPq57lmEvtknmO
zfMwB3BC86LTGVEQXYwhMVCA6OfmaypOw6NUF3J4q0Ic5aWGXaclPfKgHX10vJ1wIYoPFxfBF3TA
+FAKnMhGqPy3jPtoU0ljdnB60qD3kgZupH1WrA0ZsEvfyAXnwYwJxJ3gyOaxpAr8R+FTlDPzaN6Y
C1kqG+Lcler+D8yJoltw6Hu7u67kshJ5kJ17QSFizJ+yQ2gTs7taGWj1q8anF+zw8hoMDjrFCCoh
ydpyF8o7D70Q2Oh9z5H0A1U7/37VSZhuD5A8gygmbz4oOFAWBSzFIRR39ZPAq3z+vDIHD2I/l/c/
zuN9rkv8e1b6BZKlcoUAHRRX3lRPC5ZETeAAMRg9o0Td0dq8LVJTPlsmdGz0fx8R6TOqp1JK/Ex+
2QBjxMVlDsu5lBkt9YFrZFS+BriFbRarPum659N7bZNJbRzg38jN1O4nSKkaNbLYLU2LHPIlCA63
M5/2r3Lg0c3a30zI+L0pVEA8LCVZPgLK5d2WRWpSLVjHSL3LC7AdDgGS05IDq5vG+YVFckA7wjot
SHoBuBmik8uVkiQNQR0WOwm1/jsmFOGKSK2DBbt12yD+vxf3SCv7ORBKggqxohV2zE4hFP5mgLZ7
9fCJursASwaQjeUI7UhTNSUpYs2lh1D/Bm+icwBGQLzTNEVoLFKP08pn0DZJCiJrz1VO6GP3VM0o
4McIvwvMJYDsd2oN2kLeS1Rv3TJtesHUQQpQ7GNPXHs6m48tkiEW+6etImt3OhuN2Bmlx6lnXHa1
oanRK0iHxIJtAMrQB1yvC5o9RAPBJpSXt4ayeknK9VHwQgZJ1hFcWcF5nJZQP5l+gYJtDKTV+UGZ
JNDmPaLlqMIMNEs0zbApvTJUr4Y6QAoJB1eg8O3rgHt8yT7S/pnl+PZ99Cfwdmt093eSCdjdI4R4
Dj0F8KaJGw9qkRTBUcuMS9fREAfnO8WEHuEr/xE0cWZOjoyRN5QD44+7yL3mjbip6sM6SUVuoVk0
EZeWT64g3Zwfn9qxMktTsEYLMN6+F6JasQqd88+hEUpgootxXE1obXVy448r5GuJGqExTK+pTuxx
QwQMjpEfK2YpUTKsJuhGOEZE1N16u/pVkSmcBvSArs+cXi4izu+TqOKBYVFCP4DQvl3/PP3z5227
XOZvC0usY/IveimE7mVl6V+UNIN4c/DFymiFPrszkRgNutlz+X9xaF/o/kFzavExj2YkFQ/06Uzg
6J6ceAeBy1vEZLNyHinsEEmTuxDmwbMpSJQwdckqE9iUeHTRdrCEuRu7swL1LGrpOWsq3/JjpbqW
Iv5yUoQY9dNtUkXCy5tKuooccNLdkFFCxPrUYkfIHfcYRhJW+kBJIoabNCzBxRNkPo5Bh8qsiYwr
baqHg2KCd+pXXNPhRxs0pQxrE+HFAV0xNAl8cCVfk7+OiHpy9bfxD6OP7czShEOqQ7+fEIAAFqez
7EFGnawDayWwsaKBPRT/7al3oJZOGPpDI96ubG8uNO7XhqOASBd5E2U/GNnwQ9zXQFwNL3tehLCs
f4/1rUT/ssoXRlvNadM2y7pD0NHRw4Fq6AslkGkPlywu4O3ztpzDN1JVuippPEkUPPjxGi3VXo1A
2jFlJSDS+RI0xfpD8RbKF8JdVIwqKPlZiU7cljxMJebEiqg4fhfwL0QUOG6CZy3qvvYh5tJ502OG
A9RyAoXCT6Tp+ETgJ/8x4zXRCpV8DaTxWIkhGICVh3xCi+eguAzcpsSRKG6H7L2SeE96ClMfxi2y
W7FfdeTKoZmGw0E+152yPLAJOCVeocwHsm6wi43yEB1mMH6W+9NLbb1PSVwqeimpjkoL9aYRkDSm
MkmKjpljAd/jKgIZna5rdDd6UtLCt/lVEPLFyQJ6s+U20/mFkU1AW55P/BbxwyBDigvv9QvHIbK5
z/D11qgGf9/+GVUyL51DyETFt9WO6+wLe26HvEWt0eBrr7NLMO69nclkfyJgpqAB/uoriuYGKQg6
kBtipXnfwGpXqsw6NDzxcE/l+LV3fSPRnmg6hzsIe0NgU0wuu35+pCSkzAjLrG6Dp12JscADAhg3
+RN1H5e1/a2cvhhzv2uB7RVWrAKrCJh7bf+yHtuNFMP3HUYN0RxuCucDA+MpzKm0ziMssR1b3J+s
h6lhi8QSkfeBjAqTJhj+a9lZVvA/2T3/FByjbfV4cbsUdw43IgOHuGITxS7V14K09BDX7YuHOxx/
XB4kSeLVMCPMtefjCzORMy4Wfhr3WTLe2TFczt/MXIUFgRe5TlB6wqNNEYIZ9voEnd8EuLzpn54K
s1eMXgJlAnRfoHDsgQP2yOQup4GkWpCOicNwQvd9GUKMYjT1d7u5COIU4yI0nWNBzkjc/nCVchef
zZyUIy6//vqYQM5iRNoXUia+G267kA+DD3s9ZAJMm5K9JtiGVuF15xGyIBYPu3uIfD+Mr0s3sh/Y
5fBUCx7azPrkZqzvwHm2TY9p2n0aZ8QNmC8+c7cgZEBuKcS7EkcQuFXkdAdSyuQnXXzBp0pkOlve
N29c+9azZHssQ4fH/7CZvyNuLd5eF0xFtMVOejx5Tw1a59gJSpzwJmtgSLvxnWm+ed/hR8yFnAKv
0shjfNYOOebtoW9JZwBxiUFmtBypdrW9t+RwMLxtQa/F+BAShzvnRRp2Rk8UOb84VZBhsWywei/h
s6ovNvI7FvgniewHKcUFDX59ttXMLIbyMagH2fG/witicfbk/Fk7Nb0p5RRfs46kylK/E5xdj1xR
zq33qlfMAxZI5pUGQstPOpVNpMedVf7PVsTsfKdcoTvgyku83kfZedoA09te59Yp+KGgd8+lhrUn
rjqo2vn+DsvM1Bzhvkm2TEqHOwybiN4iX9BLHw5fIucje6G6KrEJpZ0aFacwOUGs9xC1fKD3p5B5
gEDSrKJAwUmsZbMSKg82D7ygYklFyH5SKRdgHK8EDpUJJf0Ox603c6y/XJxq1z0FcveDDDzi9lyH
H8OZ0B5ZcqdyA88QoCghS4qXC0TCa536uzcob9fLHaARnJb8Nf6Ny+zO3TPSwoPfq/d6Le9vUEjG
X3i/40M65BZNyFrtF4f91UAxaDwRx9QpIFVBMmSGSVUdz6weUTWPgSnBZopvMzEsijgNedZOH+w0
1cPXIeQBmP23pqcFR9oTKkRzmt03RMaOo4dEO3zK8uzTyuogcdFGYbohx7QF6c+1c9GtxwAgyx9t
np9JkoicU+HoFjwK7sa+suKTATcVFbge6ZjHwrjzH5QoSChHEBLMz/bQdRwePFzLF2C4UyEDWWS+
NNpHdeAiE24X9y8hh9gp3yuTcMO9XCz+Ugxwf1D2AybfvZwE0kPrAzrMx6vfAyFNYOpbdNag+Lpz
Nnj703PX10mX+3ELbVX0+Ih6zkF5yICS+aMa/H4SIeds9E4epU1DU6g0QUBWcdQ+vpKQOeMhagqF
6iG47cK/QdiWnlbL0YzsU4GtsH1iyTyFiNp0M6SgkispBeSUuCkIcErWJqd2hUGbdjfbXOO6Ej5B
hNkzppTBusyTpS8GazHXVzlWYXhqqUv4Nazl8RE2MaBRNPfOgG9EQMNAM4hh7wD5ZBZm0uAFlsBn
fb57c1N5oI/4mpNu9HhuiB66Irmqb2VQirR+reBV4WZLVsT5J3TuxoSqX5C+yOo1d2Rt3KC8fLHH
OVTj3t9YgWk/05spWvlxIhJdKS7EilkL5fvgn+nDS39aIOeIAba3JGvNKOAUifeuU3dt0xs73XMg
wIzuulm2Uhut/61uOx9tpS19NIdIpz+6A7j7jgQwQDhzXcQxNOSOeT1qI7R1bsfccFFPxx2XsVKb
dvqUtSa7SfhaVSMCPJD2RIizwbah6pGv6aqagdQi8VNZVLXCoZ0gtkmdUSonrTOsW3PgZRV0gvVR
yBaozOxZDfvrFeTbmLsD9Q92RsnXgKLLVf3kUW+0bAHzyU3UtNCt2tUPm7Tb+N52ntNVNCKDyY/i
i0sPZesTr96hgr1W3rl4jkOJB6X5Z3XLOxO+OWcKqsZno/5tW76yGsVdipa7mzA6f9ypBNVY8ain
k1rpcefqh050p25ktyHVKC1JGVPQ9WnV01Zdo+IujGbOqmO7Q19YzYtxkfhQI4CHwmXp3gWTtL3n
Z8yIWmH5gyMA9DRLuErwJfIWgCwkfz7PpXN3gtj6eMRm4k/LcPlRxMOSvpGNs0uY9JniVhgklnc4
V4aPQ/jbuIVSFcxDyh5clPMhvTEjbfiiwwOxeymuZZ107y5NfUlXjPNWcLjWehIActyqYHu3nLfD
tU4O9K/ilzt8PojUC1wHaFFH42itljlLDEfhy1xxhVfJMQiX4bCWXwaDjQGetRXU76ArRByOKGwK
QHUeIXf0rYrOIP5QF+XaCq8AqrvulDv4IFYHT+EoSdRw6Uhd6e9XARJRY2jz+Djdg29Weo8FtSpN
bUUnDH+IXjAek95mg1VtJgxvdYCavVdNPhFcw2dd3/IHSasRDCoRWuUysfBSbLRqKiE+vykJZbJf
SS2JB5u1N7GnWCxRyg5OatIsgl+NXH1B4HV6Knv66/sYLjJ18ASSHTF0z/SF2KTU2AapM68u2Jv4
70SPStw+BSE1XgPO2iRq7xiHpgONXapZjSLEg/cb8iFZGVRhoqAz0SMA9S3+eAAL975DwW0xgnMv
4vIRdEIOfPI3u3wfHl2LggAcgfMwaJr63z5l0Wlk0GpEl46+JLTjcXBp0Z857anVPE/QzHRjbQ1E
xdogLWs3NlXge7LwUBgea8wjbYUnkQTBepdzNwA5UIVIBFUYtqg7BdqvkhHOXnz/MDQMpRTk4AZw
2w8WjOKweS6BeJsOSBiybBsBCG41auAIb7YBjcuQIzacwX1madfdIAKXfxLcIifdRwpNfxeNBU+F
XyUAk3ravqPnkuJD6c1smN+P1sy6Ftw7sAYEylR+gld6qFZejj0gtZRbMlFFUMuiLjpAQaJWddp1
2tuyojasxerEloxJAQxY+P5KV4Jb3nZpMsiLf1rhQUf/6S/k1g73YbWGe/2xMsUbgb5fYUNWG6FJ
YI3JJuaT/V7Buu7bMoqM2bwFyYkcFA2I5CXt7stlWrSRLRlNt9Pa9qK+PhBgrmtMB+pZODrSKqxV
d35IxWcRHbUjUUTUQe80iy7jflz8BMBdInJO+rWdEy3uLlzXAMdwmp+6HQZm2oQoUrtn5kraU3V0
0zRGOZuznhbipc94YvYICONh/Vy62XmztSvx6mBscQvKZH/R8MBLjdyUyoWhU8DK/GQyomBsvUNG
3SeRu1jUEB3Z5tO9sSgbFhcJI0DdI8S9AgN6FvBer8/1a+hIVK6D/SnAqV33wxlM04mvdXlB44nz
kBfZwyRnswBJkXiQc63uyGo/V29TOOygVr33PhQN2lWUcOMOB/T66xfCwbdtFytl4NnttlGF8q3c
HClrrlkxbQvEOcle+CrD4yGjftnnrmyMrEu9vlSvfEd28RdY1FTdo6/7PQJYFxu1EQ1vfGg0MbE1
rcvg7GnhT9CpOFBUDJJamjiSWrpW0HjXluVzzLipLGQlyWT8Ei14MXCBC4OnnuxuP1jeWMIuYT7n
N8Q3hNzbqh8utl/IjxrBGeFhw5gOA9m1TMBdDdhw96DlY+jva8XpICDjz1Dcw1QUqt3HZy6MOleU
TdhrVe8dzPcsPiyI/kMCUD0kIkFQpqsPwVyzozQQn1GfVS0+D+gU4DN7znN2KyqEX0H6urD9aEQW
NLTIaAcowYp/jA0iNVGSGoJ15lu00a+tpj4xBPhcMkK9DAss69fuDrp/PEbMySOgd4nnmUbFCoK5
vPUm8EwP1Votk6FQFfX2rPMw2xogCvraGOHaH3lM0+Xe+L9hYGNnwpzCkIKc9yYA2NFJ5azkdc8T
XcfU4z74ezqRiVAu9AcdbvJzhzABIRNp5zwKIPhmbCjEbMmMdFGUH4QNQuhQpCc98FtU0NvG5T4I
QZ7gfeNJ9Ao+3AHYke8AP8lkYKjwRs4MpMJjVlkhl5jj3tP8t6xOMdRnc7KI9T0NW1065DXPa2DD
lcVIpNFS5w2opnrb2hiJAEbo2b0VhWGwN/gRw0xtqwC1lGspT4gRxUeXVvBYydZ7LlsljbaYpRFe
D8jZryRGQq55LJHY/s1Mc4yL5TeybHcvOBVTy0yabpuiKE8mrO55EBTeDhgLntaXlmvjK77fGqj5
/FBEbruKN+lAo6GMG9+pxrU2hF5fGkPqc0lJy+QZZjky57WChO2TRNkn8IJUsfVZlkOUn3cNkjQW
BXavjIGhV8pAju8LEuIwMxnlIWidVpFcFFLV4/eNCx+6sMGBhpL76ozW0Cg4odI6lWWNbmVdTQ5O
TisCPjfWNz0x1gj9pGugV3Sh3sYXX6Cx7qW7Wa5eRtAIolLq/0DU/T8SjyZwP2c5XBwu/UFpDL5N
d+JnxXhNAgjoUv2dGltcVap8WDd75xYlTUFU20sNdPYUGwvqidtT6gNwo9jRet5LiNngx1/DLjyg
AxJ1hEhp+bIxeIetkZoYHlBHbQ6ideE/TQyH/Kqdt8LAYMnInHRmaY3yFzonamuHnZpoP8J7dhBf
WhaDd+eMA5wxWPpR7FKUyYy19EwatpRXe3itUx1gk//VvFHsMavQWwXe2CPRxWs6dUNg/AFy0EYq
HWrxh3mc5MzXT/TFXzVqW8yFUXNs1ZIENgun7gniAoG4KHUyMYfv1YjMxsVtZ+ei6oLAAWAKZ1kU
0mqPqUTZtvV3F8Exq3JKJrThM70AqGI962pGRfh67xF3Bs3e+qQTrR/XWi4PrJ93hzet/SZWfVIy
gI9RpRBPfjXB3Ufvu4DOPvM9DIBHK8WvftG//s9MadwZrYnvZ5E9R8OaSBs/fDG91vXEQdGX+Hft
AdXZBYFyr+gxUNOcU3rgxsLgxPtuUG31fdQTN1uTSgpKlm3N5qUBUfmRihJM1cb9H/rW24/8ayEM
plPkBwFlhfdfW3vCZWrZ7n7fheqed+rRLola9uApAhrAv/4O5KGSIteBc/JvaoZjjkDHybjay+DA
NiQ/NsASatvT+61kdFM1pL21nz3IG7/L1WsFho8FL0HTNFL/AmbmMOmOtIQJGqkIeVHsF0rYz7Qw
vy4wmw2CwSauBmPfJAMstPBL2TBo80CVEPcDq5/68iLmnP1vf8HMCV7d9CctKYDtdTDx5N1C2xjZ
zzQdFgGcRoHCad4qdXdNCMQ7yM7fryY+57ljJXSBNKT2+tW4GdubUVopmuG/3BhD1vP4WxoJNoMX
ve/nhPG1XDllJMLn7CIB46pFmsIbOGIuC2pBWmtQE/G2YNmeSL0sTgyvXtqiQ1z/jJicAuT9mT4p
n3TIb3U80ugcKSJBv8ID2egTuXO2h9fsRhxDZ26ZX4qiwKsxKPyrlgWf915S+VUhlzQe5lT8rU/x
439Zz8Vwj17+pztZaLt/KWMuXx1RhuON6vGsrnHeTAntuUJCGDCndF7FDvwul43/IjaV2Vt/gL2L
vH9ToK4muDQd74DOqJrcWDs/bV17Vu0BJvO9lPrW0zOWTM9KWaOOsqVr/q3Z2lVts0qUA8ggEfQ7
HV7I5HmLZMKuhvUm/2QxiV6FDSnlLFpn0KpEZWEnFrUujmMiaAHS4lMA2UcuyQBD60uMxsZvA1S4
+QnWQpOyjei8sKuV2H5yFYQ8/2S2d0shrsBO+72WJACrMQR/BYkgAu0wDP6PVaUUWIQNDoAuFd/S
CCDdQ54jpMEhyNk9Hevmi0C7MXPPAp/nVf3zT5sVTfiBEm0uWAtVRRIY/oXyD/Z2cRN9ehLCTCSU
kHYa9MfbUXovGizJpYFqWdnO+lpOKo5X8M9F2rhU6X8WLqtVKqRrJ7QHBBUZ9JzhZ0cr5etrete5
B8stw3P/NdRSz49yVYnaX7dqBj0nvQo3cXzFpXGzIqQ3HFZDyqKTzVzSvev48d9wwH9fO2EXOCeK
pgng22iFTwqxxMHX1oFrBuQhMk4f+KcBnViTD4cQu9sevavEJrbesY81RC3ls8z+ksL7vLTRnezt
DjfcPzXdfB/+RW2UqH5NAGO87c9TwQeiE7UpGtRLDX4PrWLumVyt+I4Idjh9kt/9hRox3UHSG+un
voOkfJCxuE1jSVkOlHOHLeZ2qmi23tjMNzRi54/3aHhZSaZGsBs8fXZvJnjLNzVN5wVz15+BQ7/U
uGKAegvUkXp/1ojZQk5YlJ78dzd5xplqgiNj4zlWAhzyGbW31aHX1v5Rk7KEv17j9hbQPYAN7Uun
wXEp7u6zRS30nwtkRXivT/CEshIPCK9pYAWzuboYGQ8Rcam8C1AJ4eYMOtva7FuKZFq0A9DGJFq0
+NIIvooRyzGS1IY3jmqk79u0dJ3cdoZGwnhKw6qY2QC1N5CzUk2UFxc17PgALdI7lzHrbilLPc3M
uqMpt02CMXNm+YCxkrIaTM/w1h1qrGnuiqqqny11O/8zNZuSuflnR5WRI+/11LB1NYpqoCj3brI1
SsgODbGi7AbSJLFkHYxSOLdVjB1F7sVHSwpKaXKGqdsWz/Yf8GpDNc955LIn0mSTiCdJ4Say1Id7
lMm5jq0RhaYLZoc+EFB8bKCbRS+rhRiYLqW+H2e8m1lggefnCSk17X1X909NYpNUxErvAXEmEUs0
vjonWgbQNNqp8mBZrPxGuYJw9yJqDZytKjiz9H8ayDz4zQBurNH2vh1YntsBAtpPZy4SvuA3L0jL
8TaMafw3H71w0noP4oZsdJwduDTAuptNZWbfiE3KbrVDwTUlRPXiuufFzS3PH7WfM9IJrfeafDql
7QmFSMBcUzI3ExYRMeFnUuXWUxCneDKAFyYN+FBqswImo03ht9kG0ta+Y2nB9+WAsl7eO+18ZZhg
doD8eiKarnBh1cqehyhhqzDx5mJZtFsc+/dItDkgH3ealk5ssv/axCfbQlD0G0OdAKdJOcuBmNJ3
FPL2daeIp6UWpkvQMVIrAUZ6D1VIZIu/9niWdDQvgtW6ZfI218dT5MMkYBq4CgroiB4R3IVZW1wD
L1jxA5UvMCzuYwAB3Xc3PIgDPC1hWSUciDptbtxBHF6DYig1EyUwSMYdfWtbkBwoJk/6QSBp5ak2
Ly46ho2f+Bo18MlkYUsvTvgH6nFzW2kUN0gIOvQTUjhxX2UYYGBGBU9Dnd/ce/ih2QY+0FuAeb3B
8omWFYnJvtfS8vbOCSilstmjZlsQkclGJXGeonVwLyEuu+vH7dpGFFaB1Vrj7QtEUaPdVaynrnFp
DsS6oK7s8xt2+knc/bYL4uqi73l9DgxBPaZGnvxsqfMpYTWWnqdK6rIhfoKwKVUndfpUJKUL+Grx
TJoEb5Tg2EK7Z1lM740uIKTplos6kqcizzCWTYLaiw3wmnjHFTGe0nVB6Xo4J54Fh2JICnJ/uhll
Fwqf5bjdoheZsAf3Cj/JLqfh5SsTVqf9MQ8AM95UZ8LKQ36bg3u1w0F8eXYY3dHMP1FUQVxnUUFb
DCVOG8uPuDsmC+++MjR1XRwKN+3aA/SbLsCTfzkmD0gpSlDFv+x6FWUP1+vHUUNdb5cvjAG5IRu4
OZV6IxrZ07X4DJkraFaIUhNx+U9KF+DT5z5UBr9VOX3u3dhSFDWunrNiWigJ+XD9/9EzwTOj8mMh
3OQXrjUyoW5Nawl0xrSo+O5KEYfy+g6UizHVaJFVNDGtuzMtopmR6ZyDDtG33sRMaVMRee+iCkO5
0hiw46koRebtTfcgnAlOt3TYmcBxHR4Dt1dOlS5wrpfxU8jITnqmHhRUPgGOBdU0p3DUWwT4flzq
r8rNqHaGobNw7L9o/upCrqlLsZXwx4iz4WM5rH5tCVp9L/KQ/i0mwdW4njRviy5RwYV6vV2FwcEV
2dS3jYDci/cXQFEO9u/HJrN/dLJ9ZoIbXpFfjwSnJ2lNWFnicrT9s4PKTu3HO8IyPOwOgtn5itsG
wNn4NWWDJV5qF2FNpZqNR+NIV2MiC5jjcBNchG8LtVY0c0/QAMoZDViB7qMkKu7hQfNGooyNQe0H
dlJAB66OeSJs1Cs9bxgHmK0U/tslhMphiHk1Xa9QeELIMte0qZBwYjpF1IgeIVU3IL2TQO1fG92I
JOEFPLZ2HlPnfuTlGxoyH/uEpyXHv6chC37XIMthXTQXNXlxcPRqcRBTqt+LtHyNfSmhA7Yye7AL
7+KlEQHLt2aEb41jO1OkEN4+UI55SjBAMYG+bKN0yExy/9GDESXywY38ufwmIGIBJkWxWHNpu0g+
PQD3thcRlCiUW2itqzmWWuzHdlEs3IublRZANkzyjrUzKOTNMZ4PQh0TTdoz+0Kg2YJGoXF0AuYp
bvqdp2XCPnsumCDhS8sfVWIPaSXIRo37Z2A14lPm8HUE2LkBA+ZOlxH+aX1r7M53BZ6HI0oaw131
2LSU14KHrwCEOX5DADPfIHN+i9HMWr17/eg4pBpEOw4QngSpx0HZv8jHOda7exX5+tFl4GYoHuOm
ghLRemxHEL587+5HleaRHEcpccK+PJhhX6z5r/gSMY299vrbM9NcuJMtRS3evh3WPvpVMq3Ds0Ch
JCayo6g35hIERevEZgA4F3D6aANCTwsJsG4UMjSUtFrmHzmQE3c5WdUkM2EK1b78w67YahL9nDNd
NJosKfQ+mU9dDFebM16inHieg5VazioAoNYgdfBnWp0PbWw0z93v+3py/4QM+4Spu8DZItvnwsVx
23MlQwQgDbG+Ywp69Y4ssS43e3A/u1Y9DD+aDHVqKAIoB+l6pXilvGM+ASUMwoNBxGBC3vB4b+Kw
Dgcas3NloWO97LC8i7mAXS5TWg6ii4RUP9e8lY8cdCBJOJcujeXCyE2aHsY4b1Njg/q+6oo61DT1
SUm6Eqz2N8N0gyk47600GHJv9Lmo6kb6xzE3aFBVMA1n815rVsT7LOPYPruUVldClZzAF/r9XDIq
5Q7bEpFdNBnxLieb+SAC1fPvBDnIpJ9GgBF/ANKJMNL86QMx5+Gb6Fr8KiU3i8qBYYxMLzBmUYbM
SWHFs+o4rSh/r3AZN7RwWYxUozb1oV3lMKtxuGbKaHGP0CeeTKNSPNfRhoGTLjZ28p9QKdk2j0+h
sSA33bIcZ3kBInm0nl8KFnNrVEUZ4WxaUvGLW534qdeZIX0gsKwi04wQGxjvkw3DOHjp+Y4B+Cgk
EB0bARnqeqU1TEFkN2UmZPvxCvu4tYIFTqI7V9meTmqEi/3TVNBlFwGp1SiPrqnL16dO1m/aX7LN
LXL7l/NgctAzjszmrb4A8wGCC3TQ26yaiQdHCU04xxtRgCLq6l7wU/IWPn1w608B502xNgSEeuV5
uU6RcHC62gedNcyRGFbE+tNf/fOdpe69Wt6Gp49D8KRsYnrEJQh7h6WN1U76Sqa6I+pAw8j8n+9o
kH1M4+zsLCmkUjbjQEFZkYdyBYU86t314s51hXchWLB4o4wB1vHkP6A61zOdVyGOjjesKO0RP1jQ
S9V+nIM5o2hYBd22OeCWyXKUN54n+nidEziQy0qVzl+s1XBEw8pUud9l0i0M9GrA1rpda1Ah4eYo
EfZ3IPeYGOdUdEVVrep0RuWUAquasRJIyErJYC7ryXo4rDVDfIaA320aSlyAOvmk+yAoAkiPfqEs
4+Sw2FbEV7MBkbTaJ4VuAbjIVdpT5R28EHEvj1OK7dt+vaAPAEYp+MzXlUsxkUTR+YqoXYwBG7Cq
ismA3QeLkSh0+ubxoIZJdf5lGALowV9YOAvZqPf33e4H7u393U8W/MSmpJyyeBV2e5jcRqQv8AV4
NiWlPQapOWFp7BqJxyzlYHS2ri4D87Te+P3vy1L3xTPhyzOznQoTAncT5k3eaxuBhRM5hIZ9oP+u
UHTrJ64lftcb1xnVb8r8bi506tveTuBvTpxjrCfz/VwDuBqihieW25zPuPvoRgsLPY/KpFXPxAeQ
3oeBCbtYcvUsEhlGWkeNbq5x6r0vUN4NOYxDzvSibh4GeUGp6Qa8iAB4RuVTUH99oHPhJ9fR/0fk
np0rohu17YHQ/0cNxUAdvc8sBhmZhEkWiVAa6bbxM3lzrPOKYE3ZbVvRJVFsZnHB/iFoj2a0zj1K
QNzGnWciP65yVAxvQQrT98dQufXwOtva/RgBhQutdJKJX3o6JT+07QvnyWG3OwGfBy5JnLT6dtsX
uLkE5FKvwA8Wka5iBezvLLbdldbwv2Cl+gSRUWeRIPiqyyjDAbSFHPIRtcZqgBgyH/FvGExzS/oH
IWc8WUQpVaOZfdYC7iEboeRSJVXYsX5tCpr2UWxOsQyUrkb8cK583hAKVgvwn6t89uXK0vGKg7MF
gEmC0iyHjwVpw+a4zPBsW1tZM9cF0cnEoKB3FmP3sWCcYOOwsAA9rgLey/gErCRDJ0szwvoWEZtd
DotwrPkheOoREXH+ybjqlkuwasdIulx7ELkdM1j8mC0HD4WGlOlJbz7AkrmujOQItoWbjhXS6HdR
X2uISXf4QVpzOfkPf5ax2c+sSoo2637ncLNWytBfMsAZTq9n/cXS1V4chjYVIRrXo5Gb3yPc4lLO
/9pyqkgFEkj0F67/S4QluFZfT4o5ZNz19Cs76AbRcr9t4mw8LALMIFeVyFAnvRSJn68ciGBxyQRx
PPCwtEHdI6z1FTx2VCYIn7Dt7K6CMqQ8jExotXcy0CioouY+se/GCr0qzEkib55OSNH2lwrQj1j7
4srpSmix6EChV2q/+p8knzAx661XNQ5V7t8PcFZ8CNtfcKF5nXmiRowrPE3JVmMOj73t/QvPPiKd
I/tP87yfjCicSZb+a4NMIWvHh56dhGux29U7FGOQ6MzQWQA2URbNisVpEAfa+8RWJzCZnFncseRN
hXrqeobevZD2+wEOE3pljQiDFDo287CKMRWZb8gL0yiHb1LF87JpftclFgYdXwl9WBgmCMTgwl8M
pmLLgyyYwOzK8yM84gQrAQ/PFiPMMpv/eZNAoDvLInMPE8Ki/DDlMNLWW2yXpM9N0eptwZFqVzax
HYJL+QB3UKTl/f4AEtEv26f1UMBC7ESbLBeci1vAYF16kKEhAW3n8eF4QltK0a3uyNnHC+OSvAXU
BYDhOU25iNOqZ99uXWqRDPfYIFmQZk12/EfeZjhGh6ZMM3Ug0r+LytqoORDiz/e24zgdyzfRfPJe
x9Wyvl75JtNL2FEUPGoq3m6DW88fwgobTbjRynChbpDvYBaI/31/CBHCVOAKZlJevVsoFeoM05js
GuRcgrEq6up8eqjLcHou71ocjt2hLcKWdkw9hlv2aIzB37pWomxy2vWsqTZrBPMX5xlwSXGFcunA
pFWAK0w3nzDsMWvPbzDSXtIEmB01yhgz6HiHHWvv99ZaOzsfpfXtcGuzCaDIjgiK68q2hiIrcTlC
YCutl2pDzi2YwC4vG2GwDBMCKzzhR27JXv49/1gqZCGGdbsGa3AgISApxb0yjSJ03Y4Wlej2T2Px
Dgwvu7y+GJL/w/klqsHuN4pUCtCW8iwzJXhYTo/3BM/IvFB+Qj18cUvbFq0Ov8AxnWULzHr+McHU
/ktP5+Vu0SArCnKxu2i796eNJO0LsEWxjC0zIopTWucmpCnSH6uizdY/oSMhc4dkRIQuttnZSHQR
1UFnXtPnLFoB5qU98nwjQcYpPdEg7JywkTRZGqre3C7BM/uhtMh5ebf0sRBcWontGXzNkLf0jrSl
RjN6PTfL3FVW8dZuCzNk7CuTf5s+Yg+mPGguB397Ays4Bn3Q4Cz8cY10YIeJPs8hxBeKAhARuISI
IR6DxQ0tY9hB7PV00RnRld/CFVeME71rJtafs+c+IBVagFEOcdXJKP7PF34DXR8zvCMI6GyC2DjP
q2Bb6jR/bpzFPwT4qfob+o/UEyzCgn7Yd4qTIVFt70qRpFOci93/QCxuwKHMAua5EycGTiae7FL/
uj8QrXvJj43pkUHpB79bpbrAu5dYkBOYBseo6cexSWm7HRKWWh7XA6Pvcu4MpoAdgbwABEa05C5D
HH0rVTXj7I+eeIpdGPHs3LqJ+wLLHBiCDRL7qriC0Bqp9h9zgE94TupmUIU4kjSttx8y0KjFHcN7
vTA7VdspUGKgmNiZ6KvkMtdd6EweacXMz6Fw+5hIIhGxWS4d6+qI8mfNDZtNuxs9al9v6TjvcI4y
0TjNJKWU3lnzHNPlfFJ0R47NF9oACnkrqvtWbfKM5nuwwZAKhnHYIliqeniHkEVn2fiDhJW9ARU8
fh/M88JQnpFULyLQqXFundxspMjkCKBDTBZo/98kMfRIOfrFbIFiY7ZhU9UlS2HSouAJmvELEXQ8
bcoeV3b9d1GNoUGW0lF8I9lLjj1bdXg9C9+2WazFWHf1HFKkiSMTtbkU2zZjaDuF9ZPQp8kAEcfW
9sBWrgFcC01PjvQspW3duf0Kt+g4Hvvxo2Glo/pSZQEXMuCGhElCV28Ucmj3nOLUwS5OyBxuwDcz
FKoCR+mJzxaOb3vKP7AVvBKJ41mc+qwiOiVPKNmr7hNJCZ18pBbs+Cddh/kLsIEKZgA2jtD47pSZ
p5KCq94ZDPyw3Nop2I00pBsM92A+MGsnQ8YEBr1YFkxhCBt+57FJZEs6pvVc0TKHb1TJ1t5N3nXr
OX6IP1JZv32lvFmijCB96nEI6Ou4IXJVTH6e3qjBSs5NtJw/flVynxkmHTCM1yCJhw5SxCEfoGSQ
vqjd5YzB+9Z+z9lt9eHlqIooTwc+vSNLzu2C+JQ764wW5uAIoy6hnXXrtan/j2C7qnx8cyAN97Ad
6IstGCUlZ6EJ764zJ8p0TBCjDxMARoGF+3BUIXlkYvnQvSRTAg1SB5BgTE1VaWNmfus5kGLL+3nm
d7GJeQ6Q4BOzDbLU9QAEi5V5dmopb7Ch4fvaYL5UJVMo8q2Wd5T5ktHRYCT6Kq12ZGV6pe/8zklw
nLqzmcTbXYGzEzPHehw5qDqHaBJJ/9bDanCCaVRwmJX4xedzmVIjWVWA4hr/e4poW8aT5YFh2xMF
SadykJUpdfVyTsdOGgdDZ9QHv8EyI0MpYtsRoiihEAADrYmosp9aEoHj5mEIP8KHFh82BMwc3ras
ZR5VNJsLweQbTaa1nlxPIze4B1y8jnyS+uuSMxkepQPGdBTYEtggWoF5ax5KrUjPMr8CRXGyswis
5cBemXndrXcMPxCRjTaME8ZpoJXBvqq6tav4MfezuvYIph3xEbwO+WDr2Txzrkdxdx8MahclhEKK
fRmScWwQLsEp0P8eA3NP6QVl62zHccoENknuxqTG0XeUi3iMgnDz1d2t7qpj32zrHp5tqnEpUq2g
+PrY89AmZ3XJz4VuVMOZSPJYc6mjugeyRasBWRJfYY8QGpzgtGpNlp6EHz8HK4Am7TnEY8bRZoLg
XwSBvj7P6CXuhIMasqIH2BvrI6CS0fAJvH3Tfr1JRdtGeH4ie5SoSozHDP6c/wzfAksyZ9+7J69x
iJnRXWXpxlZCIfB6ACoLj9Nw5g6BvFnVOOJ1D7wiw1CxaSi7BNbwEvjZJsRfm8w53QjT8XERbXVa
fB4wdXM3EBAGVpatz6Z/abFERJ87CFgiEIey/UyfOvmO0X2dDZglv28iNf0WX921TnHyvGFfcVSi
pto/FhZlSnlvP7aq7lJ2+ivqXAJF+FNGrYQTN93b97UlORU3MsiAWJ++2phxMN3/WrO7aW+TNa04
DzGuZ7wqZNqsai1/6B9mPTDGeD+yUwrMvtWm4nKrsN1+g2Sh7dqhiiBc/Wnu9SLbT7zcEW7SVXHI
mt0x6eYMIrs+wMeFlNQQSEQyuDnyUE+Wfdbu4yucNVx0UR4O/eAeQYLrfbt5uvizOIKdpyy0lVNx
LLj+wbdUWNB4zbftM8qZKWpeyz9QqZ+7eEZz9w1G274/vmGLqcqu/5VDhYvRZil3lcPqnw8qbgYX
aXe801ZeWVc6WKWu2nmVD9eS8hsTq14fG2A+h1RM4YOxoMssq2DpEGTpGqegc09W2EbVHtyd5Fqt
gpwrQCmtN0alGtTiGkBPqMBsqw+zp4tb531Rilh3KnrT4kVNRGNtyCAU6NV1yjuUXjCxU8Gzvouj
RVOawtqPTCmn4s2229eCoXFy2kazJ4yH0gHLgP2nAO7tmazj6pnlsio/viZKLyM2Rxc4jzKT3zw7
Iv9mTxAJkvgIhF8Hx8E9sY1D5Rg2zGza6SRA4W1kpY2z46JruGmYDvmwsEVRJ8PoPAQGysqxrD5R
RbV5+vyuabise6KNoapyE1xJNNkIdxzDms88Ufr81sI/t1LeA0xSScaiizJBF4Fwfr8QfpmKslBw
DXTNLKUDObjS1PUVnSuBC/cF6B6qoHhy73llyxB0hflJ3FCQ/t3vapxdU5jsukWXdtSuitDLSJQe
C2BR8yIgm3FI3b2f41Cq7IW0TFK/7EKdor+/cNMiqdT01wSJwgXRSvxxhJnxZ1dA+QDMJwrqdDSH
QjLjmCP0Ic8r4UoviPpb3mUo8qPm75RM6erLTrzqnhz/CEkzvzDF60Pzm3tVBjMpeOzJtXalcWS7
nFNJEkXD7XjfZF7/8lIs6gN2Mtd51TarL1aBT+6ZZUdkWtfaUFh7v3Al383TareSdrWFvn5OaWwt
ugr+RMCNOLgd3OReeT0tnx8sY/99y0cCCHFKKoNwdWqgj5LFJZRnRe8a4TJau0Br2/dBhwvWFwy2
hyUqhOP18glMb1yGdiM4XD0nw/3xoTX53kyrwyc1Kg8kBWSbHtu2ajAGsZaP43b+ikUQDVigR1uH
VSvKAhFA7Ntl1z2ujRUQkgFkyR3zQ+l5VrUD3td1nypU3TtQ+VnEVGIDdv2ibTk8ZnFFXhZqNO4k
gvPCFb7y2s7diVakcr/M/MurdzTG9yexU51iHEen5yQqBCY7gCCfpn9Fc26z9J7xzZOANlWEaWjA
TE/JG4bYFO5Gvoff+jL9JG5GV3T7Sc8xRcnVwIw+WX+EB4inJ8ak9vSWxcECXNz7yI9gABQ9nwM8
HY/Sj0m0kuzLG/letf4wt7572bT+paguC3eJ9sIyIWCWAraVYCQER7cPTKLW+XT9/eFswqVJGeRN
q9NBU6bG2yzjz6uFVlmU3npppiQO7m32y3g5fTDzTwIo26cadS1CCtWYzdHC10HAeCGroycB6lg+
gAbybKi0QZ0wshDeVg//YQUZSDNpwHS2n9cx995Qkq03BFws6b7+FSscFeUOSyTQUxb1qxGiwuLv
/JxOxL9rewQ4/Bdk7zPfzqkU1/Rr7Pzl4L6cDvWQBibx6lQmwu2LIMwn94n7NHGIfrN3kzEslmeP
7MR9BbZ7sTMYER7Tw4ileC2HpcxknipF57US4SBbo9e4+Wb7olWkp3qeoyK2angPFXZxgbjptPUg
7qHxI5ZEuLAIkrl5ay7Ko9jv1h+9n4Q6v+9k9uIE69arGd7dnU6Ktt8Q9mplW37T7G3aXPmNaQUk
9kJmm+lA7TZ1AgFURbwa79T25djrShmMpNy+Fc4ut3blAikQ29aQcXSh7/6GAeAgdeCJO3ZTBKhf
3jrOCU00kPkuF8mWQpNFaZ1NICi7pwxzfe/8fO9ex8/OW+v2Fr6Bjw0neZNwRkpVXlt8tHmMPEBB
C8mCMwW3dLOV8M97fphpqLDhLXDOfRa5iycF/Pp2KDRQJqqu/IQc57951KEoiiJXO5UAKseBttAE
W+KCwC1P2J10Y5wPEa5k2fjhQ4q7G2WehYMHa4p4MNa7gcI6nDWvIVuR3Hp5A9o4e+lqWjcXHW70
FTx9lobS3segF8y5lM2k+1FwFO/Zu1hI4q6A2ONzWHqB6+IUuhMkuPnoBWnoFAWymm7dlYufM/Yw
Ew4RfYUPRtv7CQeFr7XaW2uFnAWFaYtmmhqqhmOEmJEJn4QFA76R1q/Y4pUHZeCWq85gr5dFBl/g
1mgb1ux0JUz86FTGMhYc75LZYQ5uQ+jro/MedVoxWZm7jBGuPYZ6vakeob3nhQO0M/WhVXOVZt1h
H7ZzNFfBZFYNngmXFgIEpYcaebC4d/ilR0ALeq4FoPqJ+Hg/XG+yf8C2CBxYkHOMHNSSC8NoTEtF
SjwDmmhinIRkuIDbomDljLzG/2Wm/HjvRxDpnVzKXBxTNXQku/yDXxDQHAbg3kR9lT8n/4PJHobc
uRaN6SkmXAcF3airhb4CJ9Ncd6tcgXZM2kiPMEdN7+rCUaMSo5lim0bDewhovf+lI2aeLVdMo31x
J1wlMp2b47Xf6oL/eo6mTwAdpc2HSK1OeZjH14od6HAU5ZROoVmhFxCbSXGOKGYzQTq6HcHdbseg
+nm6meHIkq/Y9M1UoTi0VXfbPpOAYckvamuZi7pgpKPa75rjf5AoE/Jd4blkDPwc/wYiE7EtWG0y
V0e0nEpDZuK4e7iBHwpeaaGA7dQBjcT9jLD4f5V9P0HhtZxqM0lC13UXEZsLqu6j95hHqhmBSIOv
X2W1Ndd6Kt/oZFrMdA99mnNo11k9Iue29DK5xGXe8KBdae6VzNOZVkn73wa6uRCPqjDzhn1xVICV
peSCgF9o1zOWr8UUTAAXwNkjYZI+khvoYqE0DZCNni3JORAKSKTJXaPA7ms9gJzI2y5Byvy0Drgd
A9g+hBbXGQGWlXVR1MKMxa9OvNRhs4RzWws6n4wt0xEbdev1Qh3jKy/2LoijwgG2ftUi4kFWuyyS
nuamvY8WYWp6sLxrt1yVpkfXnWvQTv/hKAxDJSDeQCRgT+JB2AJA0vLF+7DoTDdt4iL3s3NfcQqD
A+Mw3FaDJzNpBXfpumtqv0P3L0YGHBjO7duZPHh8dElxsdbPylsOLV2XOkH0VWqQZ+oEz8MnEISn
SKBbaN8uYyKwJrH/J9oTQlnMyu7bqDJ/87nH+JmcvZ67pnDvSMf1Q4BEDGMQWovaTxnEvqZ7YkjA
dU5XQtlhMBjiodRBNIUED7Mqkucw8+me28fA/a/dW2ZfNpyXcdkK6TH/SV90zQsodJRsff9MxKxE
0BDB2izzj3/IS3w58Vz2oQtODofUX5a9WauUa2Uzv2EAopiVMlrMSSzEPEVhV4WZyYMFuDiFcO9F
u4ZHZx3BSy3IAt7g0lFhLOCcWDDhM9lCR9aBp7sEJUyKL3vp0tC7oSpuZW6PEkUlx2d2eAo5uLW8
++SBe2vafgZh/GOTQyh3+9URzvbs4NHy3bvKlldZU0NphVKF8xGDzuHxxpTdW2RRu7cIfqgDII/F
3Zyp4I2S6IHUH7wPScT0cFiHgbM36bCBK77TdAQe+DoD5so23q/yxVcBGGO/A8+1FJnjyn9ExFzd
OqWaWca8ETtg4AzXEsZfmR+LyuZg5JPTxhyZ3STESTUeTyR3eKzwsQJQV3GNlxUeFhp6VcDSt649
jzkHGekAbTB2GZsqzTu+LcmWsCY/mqWCjPf2022otB5v/YZvru889gYVCrhk7aU0+ZLds8pFpSDk
JDzGX+lc498iEDJ/VPkn8b9r2QZXXYTvvx1Q3CCchaXIDgq95ERvBz8+bnTcMl4DnuFWSoKRqXPj
vsrnCUrnuD3OBJ/uBbzXEEsyahPHdGLzoJGcINsXFfKom9nMh5s9Df+XxCk5puA80S6JTA//wkUw
bLyoVwu6EN9htexi2+DzdbR3mROR+BMM6tRqKN0oWygQigQO9T0EAXF4x1YMfgg7slhHma+DpjpW
AedHPVvrN3I4ll8hLnQtLpZTCWaf0nGgHQVU7rRUKocVER7NCr0NRILptRw0fGB2pXX9vMZfYKnc
jbEQnMwskUMTsOkjJnH6U1zOF+uT0AjureNR3Q4SlnR80Bfa7jVFmag3F2CNxHMZfN4pZIMDImMn
rtpaAk46v+5+tXkmf+2XQ5kBEJWjQxPiLPq5bIFijQwwDAG2RW2crEkisM9pQ7UErCfS4VGozTwI
zDHMgMvUKsHgsKq1eNcIO6XjfMa6KMss7m5czF4zksVseUuPDqifqKce1x26Vd+pd4zHZvHpprYj
DEct0cBV/GrLxa4qjmisu4vnd3pVNneV4xZkz5wguWAf639DK69bU572ms3AYTp4Tj1RwxjCGAAq
ww0nQIEgPqQpOOFy722MYmk8oe7gU5pl9dzJwkSmxQMwCUcL232eWyKFvMHBvW7m/gsANpp77TtE
Uv1xfKV9DAZBKOUCuskk5XiMrVkg1YjD5kgUTbTzXs4wxF+Qb7skJNtAJ1VJVbPIpT8CZiFb4EXE
8p8xefzRFpi8sxcE4RFg+RDgievDkDlCeBRxdnmzhXSO/TT2i0faAQ+pyhTUi8iiq+fsVCPx7hca
R8A8YHPZLTPaivdg8n853bN9scegj4k/PEuRhcafaW2v1gBZ1ioDahcjza+XaxkHuIfmrEKiSM2w
HISPwW2zRkzuGMq57x+0VAEEDIBckNkMY7FrHS66rN9q6kewVJgRJsGwFHmaXRdrGESYEUDjGnIm
jZZ/jddVESWVmiorq0dK4xzPUhoC424kYLTkOdCrD7AZRI10NMoL9Ddpc52Hs0evuY8cKv6JzJrZ
R0JOrC9bDuFzIJhjhRE53mH2nrxH7FrMEaCvw+FKelPzKgMfPlky4tPWikHORjKeXoNiy/kFSbnm
fSz/qq9WIpDJ17KdH/8iFJMtHu9jZo8QuiwmFqD8ZXtyC/MQggRG0AVyj39/pCYu25c7UQWYGQXz
AITYF1n1fbtz6wkdqs5U3YluJ9cN3peiu+oDwsaVrk+LWsSUzSxZ/3hYMoKYVomrrEgzgWFjqvLq
KBH3Vgs5nQI7D8kc2irGrBH/JhQvBgHnOnYuG/EP+paoTPamIVxTdfQYQc5sz9ZVXoNTm9ysvOrh
k9PABXwfVeCafdvfTsSOASCfxq3ccltgYZqUAfQCM9GVdUVe7R6cY/BjKLk7ot2YpXGy3CV8Qyg1
5MBUtyuq/iAR7Tv7M1ZH1BgVZ7nxlVq/oApQ2Ul8JnYODq0zYtxFloJV2n/osWkzfm/7bBbUXY6i
IuvUzquLRJGxCEzzE5aLAwtLBf+NySF06dVW86ALHPj3S4dK1439Xhe5jBRKRKm/h87g+FoVufDE
SnGeZnMLPiXcGV5g6k+p4MeFBf5lE1Mhl2FrPOeFhuX7E0Oy1jWDBiceTZurg6cpgBCqcruvZJKh
VZvkhzubH7ZarxbX7rbUyDd1yN8jEoUjq2Z+urNP5Pjs5lWyCMIPuTsZcS+ms+Vr4PkOgt7xe8B9
Kdi9oG5kXgQ7R2f2BuNL1smbjmoxxZiixXOsQnfCXs7rlsND1GvQBsdlyaHcgdsrxJmwGtmysye8
zprEZqIkDKcUaLiUTrZathNqOBLRoKs3TF2GL+cL0LJ22NMB7h9fEypOTBXc0ZISeogs4sN72uPy
ztIrQN0rbwlb6Eer/PQwp4S1yilL0y86KhhCL0imN4UQD3KEgbAQVgV7PpJs
`protect end_protected
